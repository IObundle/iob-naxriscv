// Generator : SpinalHDL dev    git head : 6b321406cee399fddb7b5231ad722d8811ffdb94
// Component : NaxRiscvAxi4LinuxPlicClint
// Git hash  : fb12adc9d4dcd7c3d92bc31903d7cd66c77f30aa

`timescale 1ns/1ps

module NaxRiscvAxi4LinuxPlicClint (
  input  wire [31:0]   ioStartAddr,
  input  wire [31:0]   ioSize,
  input  wire [31:0]   externalResetVector,
  input  wire          clint_awvalid,
  output wire          clint_awready,
  input  wire [15:0]   clint_awaddr,
  input  wire [2:0]    clint_awprot,
  input  wire          clint_wvalid,
  output wire          clint_wready,
  input  wire [31:0]   clint_wdata,
  input  wire [3:0]    clint_wstrb,
  output wire          clint_bvalid,
  input  wire          clint_bready,
  output wire [1:0]    clint_bresp,
  input  wire          clint_arvalid,
  output wire          clint_arready,
  input  wire [15:0]   clint_araddr,
  input  wire [2:0]    clint_arprot,
  output wire          clint_rvalid,
  input  wire          clint_rready,
  output wire [31:0]   clint_rdata,
  output wire [1:0]    clint_rresp,
  input  wire          plic_awvalid,
  output wire          plic_awready,
  input  wire [21:0]   plic_awaddr,
  input  wire [2:0]    plic_awprot,
  input  wire          plic_wvalid,
  output wire          plic_wready,
  input  wire [31:0]   plic_wdata,
  input  wire [3:0]    plic_wstrb,
  output wire          plic_bvalid,
  input  wire          plic_bready,
  output wire [1:0]    plic_bresp,
  input  wire          plic_arvalid,
  output wire          plic_arready,
  input  wire [21:0]   plic_araddr,
  input  wire [2:0]    plic_arprot,
  output wire          plic_rvalid,
  input  wire          plic_rready,
  output wire [31:0]   plic_rdata,
  output wire [1:0]    plic_rresp,
  input  wire [31:0]   plicInterrupts,
  output wire          iBusAxi_arvalid,
  input  wire          iBusAxi_arready,
  output wire [31:0]   iBusAxi_araddr,
  output wire [7:0]    iBusAxi_arlen,
  output wire [2:0]    iBusAxi_arsize,
  output wire [1:0]    iBusAxi_arburst,
  output wire [2:0]    iBusAxi_arprot,
  input  wire          iBusAxi_rvalid,
  output wire          iBusAxi_rready,
  input  wire [31:0]   iBusAxi_rdata,
  input  wire [1:0]    iBusAxi_rresp,
  input  wire          iBusAxi_rlast,
  output wire          pBus_awvalid,
  input  wire          pBus_awready,
  output wire [31:0]   pBus_awaddr,
  output wire [2:0]    pBus_awprot,
  output wire          pBus_wvalid,
  input  wire          pBus_wready,
  output wire [31:0]   pBus_wdata,
  output wire [3:0]    pBus_wstrb,
  input  wire          pBus_bvalid,
  output wire          pBus_bready,
  input  wire [1:0]    pBus_bresp,
  output wire          pBus_arvalid,
  input  wire          pBus_arready,
  output wire [31:0]   pBus_araddr,
  output wire [2:0]    pBus_arprot,
  input  wire          pBus_rvalid,
  output wire          pBus_rready,
  input  wire [31:0]   pBus_rdata,
  input  wire [1:0]    pBus_rresp,
  output wire          dBusAxi_awvalid,
  input  wire          dBusAxi_awready,
  output wire [31:0]   dBusAxi_awaddr,
  output wire [0:0]    dBusAxi_awid,
  output wire [7:0]    dBusAxi_awlen,
  output wire [2:0]    dBusAxi_awsize,
  output wire [1:0]    dBusAxi_awburst,
  output wire [2:0]    dBusAxi_awprot,
  output wire          dBusAxi_wvalid,
  input  wire          dBusAxi_wready,
  output wire [31:0]   dBusAxi_wdata,
  output wire [3:0]    dBusAxi_wstrb,
  output wire          dBusAxi_wlast,
  input  wire          dBusAxi_bvalid,
  output wire          dBusAxi_bready,
  input  wire [0:0]    dBusAxi_bid,
  input  wire [1:0]    dBusAxi_bresp,
  output wire          dBusAxi_arvalid,
  input  wire          dBusAxi_arready,
  output wire [31:0]   dBusAxi_araddr,
  output wire [0:0]    dBusAxi_arid,
  output wire [7:0]    dBusAxi_arlen,
  output wire [2:0]    dBusAxi_arsize,
  output wire [1:0]    dBusAxi_arburst,
  output wire [2:0]    dBusAxi_arprot,
  input  wire          dBusAxi_rvalid,
  output wire          dBusAxi_rready,
  input  wire [31:0]   dBusAxi_rdata,
  input  wire [0:0]    dBusAxi_rid,
  input  wire [1:0]    dBusAxi_rresp,
  input  wire          dBusAxi_rlast,
  input  wire          clk,
  input  wire          reset
);
  localparam BranchPlugin_BranchCtrlEnum_B = 2'd0;
  localparam BranchPlugin_BranchCtrlEnum_JAL = 2'd1;
  localparam BranchPlugin_BranchCtrlEnum_JALR = 2'd2;
  localparam IntAluPlugin_AluCtrlEnum_ADD_SUB = 2'd0;
  localparam IntAluPlugin_AluCtrlEnum_SLT_SLTU = 2'd1;
  localparam IntAluPlugin_AluCtrlEnum_BITWISE = 2'd2;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN = 3'd0;
  localparam Lsu2Plugin_CTRL_ENUM_MMU_REDO = 3'd1;
  localparam Lsu2Plugin_CTRL_ENUM_TRAP_MMU = 3'd2;
  localparam Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD = 3'd3;
  localparam Lsu2Plugin_CTRL_ENUM_LOAD_MISS = 3'd4;
  localparam Lsu2Plugin_CTRL_ENUM_LOAD_FAILED = 3'd5;
  localparam Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS = 3'd6;
  localparam Lsu2Plugin_CTRL_ENUM_SUCCESS = 3'd7;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_BOOT = 10'd1;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_IDLE = 10'd2;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD = 10'd4;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP = 10'd8;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY = 10'd16;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_ALU = 10'd32;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION = 10'd64;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_SYNC = 10'd128;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_TRAP = 10'd256;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT = 10'd512;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_BOOT_OH_ID = 0;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID = 1;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID = 2;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID = 3;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID = 4;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID = 5;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID = 6;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID = 7;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID = 8;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID = 9;
  localparam PrivilegedPlugin_logic_fsm_enumDef_BOOT = 4'd0;
  localparam PrivilegedPlugin_logic_fsm_enumDef_IDLE = 4'd1;
  localparam PrivilegedPlugin_logic_fsm_enumDef_SETUP = 4'd2;
  localparam PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE = 4'd3;
  localparam PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE = 4'd4;
  localparam PrivilegedPlugin_logic_fsm_enumDef_EPC_READ = 4'd5;
  localparam PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ = 4'd6;
  localparam PrivilegedPlugin_logic_fsm_enumDef_XRET = 4'd7;
  localparam PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC = 4'd8;
  localparam PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP = 4'd9;
  localparam PrivilegedPlugin_logic_fsm_enumDef_TRAP = 4'd10;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT = 3'd0;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE = 3'd1;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_READ = 3'd2;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE = 3'd3;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE = 3'd4;
  localparam EnvCallPlugin_logic_flushes_enumDef_BOOT = 3'd0;
  localparam EnvCallPlugin_logic_flushes_enumDef_IDLE = 3'd1;
  localparam EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE = 3'd2;
  localparam EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH = 3'd3;
  localparam EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT = 3'd4;
  localparam EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH = 3'd5;
  localparam EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU = 3'd6;
  localparam MmuPlugin_logic_refill_enumDef_BOOT = 3'd0;
  localparam MmuPlugin_logic_refill_enumDef_IDLE = 3'd1;
  localparam MmuPlugin_logic_refill_enumDef_INIT = 3'd2;
  localparam MmuPlugin_logic_refill_enumDef_CMD_0 = 3'd3;
  localparam MmuPlugin_logic_refill_enumDef_CMD_1 = 3'd4;
  localparam MmuPlugin_logic_refill_enumDef_RSP_0 = 3'd5;
  localparam MmuPlugin_logic_refill_enumDef_RSP_1 = 3'd6;

  wire       [30:0]   plicCtrl_io_sources;
  reg                 integer_RfTranslationPlugin_logic_impl_io_rollback;
  wire                integer_RfTranslationPlugin_logic_impl_io_writes_0_valid;
  reg                 integer_RfTranslationPlugin_logic_impl_io_commits_0_valid;
  reg        [4:0]    integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_address;
  reg        [5:0]    integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_data;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_0_cmd_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_1_cmd_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_2_cmd_valid;
  reg                 integer_RfAllocationPlugin_logic_allocator_io_push_0_valid;
  reg        [5:0]    integer_RfAllocationPlugin_logic_allocator_io_push_0_payload;
  wire       [0:0]    integer_RfAllocationPlugin_logic_allocator_io_pop_mask;
  wire       [31:0]   DataCachePlugin_logic_cache_io_load_cmd_payload_virtual;
  wire       [1:0]    DataCachePlugin_logic_cache_io_load_cmd_payload_size;
  wire                DataCachePlugin_logic_cache_io_load_cmd_payload_redoOnDataHazard;
  wire                DataCachePlugin_logic_cache_io_load_cmd_payload_unlocked;
  wire                DataCachePlugin_logic_cache_io_load_cmd_payload_unique;
  wire       [31:0]   DataCachePlugin_logic_cache_io_load_translated_physical;
  wire                DataCachePlugin_logic_cache_io_load_translated_abord;
  wire       [2:0]    DataCachePlugin_logic_cache_io_load_cancels;
  wire                CommitPlugin_logic_free_lineEventStream_fifo_io_pop_ready;
  wire                CommitPlugin_logic_free_lineEventStream_fifo_io_flush;
  wire                EU0_DivPlugin_logic_div_io_cmd_valid;
  reg                 Lsu2Plugin_logic_prefetch_predictor_io_learn_valid;
  reg                 Lsu2Plugin_logic_prefetch_predictor_io_learn_payload_allocate;
  reg                 Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready;
  wire                Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_valid;
  wire                Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_payload;
  wire       [7:0]    DispatchPlugin_logic_queue_io_push_payload_slots_0_event;
  wire       [1:0]    DispatchPlugin_logic_queue_io_push_payload_slots_0_sel;
  wire       [0:0]    DispatchPlugin_logic_queue_io_push_payload_slots_0_context_staticWake;
  wire       [3:0]    DispatchPlugin_logic_queue_io_push_payload_slots_0_context_robId;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_valid;
  wire       [3:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_payload_robId;
  reg                 RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_valid;
  reg        [5:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_payload_physical;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_1_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_2_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_3_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_4_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_cmd_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_cmd_valid;
  reg        [31:0]   FetchCachePlugin_logic_banks_0_mem_spinal_port1;
  wire       [25:0]   FetchCachePlugin_logic_ways_0_mem_spinal_port1;
  wire       [32:0]   BranchContextPlugin_logic_mem_earlyBranch_spinal_port1;
  wire       [64:0]   BranchContextPlugin_logic_mem_finalBranch_spinal_port1;
  wire       [31:0]   DecoderPredictionPlugin_logic_ras_mem_stack_spinal_port0;
  reg        [48:0]   BtbPlugin_logic_mem_spinal_port1;
  reg        [1:0]    GSharePlugin_logic_mem_counter_spinal_port1;
  wire       [31:0]   Lsu2Plugin_logic_lq_mem_addressPre_spinal_port1;
  wire       [31:0]   Lsu2Plugin_logic_lq_mem_addressPre_spinal_port2;
  wire       [31:0]   Lsu2Plugin_logic_lq_mem_addressPost_spinal_port0;
  wire       [31:0]   Lsu2Plugin_logic_lq_mem_addressPost_spinal_port2;
  wire       [1:0]    Lsu2Plugin_logic_lq_mem_size_spinal_port1;
  wire       [1:0]    Lsu2Plugin_logic_lq_mem_size_spinal_port2;
  wire       [5:0]    Lsu2Plugin_logic_lq_mem_physRd_spinal_port1;
  wire       [5:0]    Lsu2Plugin_logic_lq_mem_physRd_spinal_port2;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_robId_spinal_port1;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_robId_spinal_port2;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_robId_spinal_port3;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_robIdMsb_spinal_port1;
  wire       [31:0]   Lsu2Plugin_logic_lq_mem_pc_spinal_port1;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port1;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port2;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port3;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port4;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_io_spinal_port0;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_writeRd_spinal_port1;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_writeRd_spinal_port2;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_lr_spinal_port1;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_unsigned_spinal_port1;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_unsigned_spinal_port2;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_doSpecial_spinal_port2;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_needTranslation_spinal_port1;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_spinal_port1;
  wire       [2:0]    Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_spinal_port1;
  wire       [2:0]    Lsu2Plugin_logic_lq_mem_hazardPrediction_score_spinal_port1;
  reg        [21:0]   Lsu2Plugin_logic_lq_hazardPrediction_mem_spinal_port1;
  reg        [5:0]    Lsu2Plugin_logic_lq_hitPrediction_mem_spinal_port1;
  wire       [3:0]    Lsu2Plugin_logic_sq_mem_robId_spinal_port1;
  wire       [3:0]    Lsu2Plugin_logic_sq_mem_robId_spinal_port2;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_robIdMsb_spinal_port1;
  wire       [31:0]   Lsu2Plugin_logic_sq_mem_addressPre_spinal_port1;
  wire       [31:0]   Lsu2Plugin_logic_sq_mem_addressPre_spinal_port2;
  wire       [31:0]   Lsu2Plugin_logic_sq_mem_addressPost_spinal_port0;
  wire       [31:0]   Lsu2Plugin_logic_sq_mem_addressPost_spinal_port2;
  wire       [31:0]   Lsu2Plugin_logic_sq_mem_addressPost_spinal_port3;
  wire       [1:0]    Lsu2Plugin_logic_sq_mem_size_spinal_port1;
  wire       [1:0]    Lsu2Plugin_logic_sq_mem_size_spinal_port2;
  wire       [1:0]    Lsu2Plugin_logic_sq_mem_size_spinal_port3;
  wire       [1:0]    Lsu2Plugin_logic_sq_mem_size_spinal_port4;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_io_spinal_port0;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_io_spinal_port2;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_amo_spinal_port1;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_amo_spinal_port2;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_sc_spinal_port1;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_sc_spinal_port2;
  wire       [31:0]   Lsu2Plugin_logic_sq_mem_data_spinal_port1;
  wire       [31:0]   Lsu2Plugin_logic_sq_mem_data_spinal_port2;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_needTranslation_spinal_port1;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_needTranslation_spinal_port3;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_feededOnce_spinal_port1;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_doSpecial_spinal_port2;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_doNotBypass_spinal_port1;
  wire       [3:0]    Lsu2Plugin_logic_sq_mem_lqAlloc_spinal_port1;
  wire       [44:0]   FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_spinal_port1;
  wire       [44:0]   FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_spinal_port1;
  wire       [44:0]   FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_spinal_port1;
  wire       [44:0]   FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_spinal_port1;
  wire       [24:0]   FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_spinal_port1;
  wire       [24:0]   FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_spinal_port1;
  wire       [44:0]   Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_spinal_port1;
  wire       [44:0]   Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_spinal_port1;
  wire       [44:0]   Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_spinal_port1;
  wire       [44:0]   Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_spinal_port1;
  wire       [24:0]   Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_spinal_port1;
  wire       [24:0]   Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_spinal_port1;
  wire       [31:0]   CsrRamPlugin_logic_mem_spinal_port1;
  wire       [26:0]   BranchContextPlugin_free_dispatchMem_mem_spinal_port1;
  wire       [0:0]    RobPlugin_logic_completionMem_target_spinal_port1;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_0_spinal_port0;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_0_spinal_port3;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_1_spinal_port0;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_1_spinal_port1;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_1_spinal_port3;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_2_spinal_port0;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_2_spinal_port1;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_2_spinal_port3;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_3_spinal_port0;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_3_spinal_port1;
  wire       [0:0]    RobPlugin_logic_completionMem_hits_3_spinal_port3;
  wire       [0:0]    RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_spinal_port2;
  wire       [31:0]   RobPlugin_logic_storage_PC_banks_0_spinal_port1;
  wire       [31:0]   RobPlugin_logic_storage_PC_banks_0_spinal_port2;
  wire       [31:0]   RobPlugin_logic_storage_PC_banks_0_spinal_port3;
  wire       [31:0]   RobPlugin_logic_storage_PC_banks_0_spinal_port4;
  wire       [0:0]    RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port2;
  wire       [0:0]    RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port3;
  wire       [0:0]    RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port4;
  wire       [5:0]    RobPlugin_logic_storage_PHYS_RD_banks_0_spinal_port1;
  wire       [5:0]    RobPlugin_logic_storage_PHYS_RD_banks_0_spinal_port2;
  wire       [4:0]    RobPlugin_logic_storage_ARCH_RD_banks_0_spinal_port1;
  wire       [5:0]    RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_BRANCH_SEL_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_spinal_port2;
  wire       [0:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_spinal_port2;
  wire       [23:0]   RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_spinal_port1;
  wire       [3:0]    RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_LQ_ALLOC_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_SQ_ALLOC_banks_0_spinal_port1;
  wire       [31:0]   RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_spinal_port1;
  wire       [31:0]   RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_spinal_port2;
  wire       [5:0]    RobPlugin_logic_storage_PHYS_RS_0_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_READ_RS_0_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_READ_RS_0_banks_0_spinal_port2;
  wire       [5:0]    RobPlugin_logic_storage_PHYS_RS_1_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_READ_RS_1_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_READ_RS_1_banks_0_spinal_port2;
  wire       [1:0]    RobPlugin_logic_storage_BRANCH_ID_banks_0_spinal_port1;
  wire       [3:0]    RobPlugin_logic_storage_LSU_ID_banks_0_spinal_port1;
  wire       [0:0]    RobPlugin_logic_storage_ROB_MSB_banks_0_spinal_port1;
  wire                clintCtrl_io_bus_aw_ready;
  wire                clintCtrl_io_bus_w_ready;
  wire                clintCtrl_io_bus_b_valid;
  wire       [1:0]    clintCtrl_io_bus_b_payload_resp;
  wire                clintCtrl_io_bus_ar_ready;
  wire                clintCtrl_io_bus_r_valid;
  wire       [31:0]   clintCtrl_io_bus_r_payload_data;
  wire       [1:0]    clintCtrl_io_bus_r_payload_resp;
  wire       [0:0]    clintCtrl_io_timerInterrupt;
  wire       [0:0]    clintCtrl_io_softwareInterrupt;
  wire       [63:0]   clintCtrl_io_time;
  wire                plicCtrl_io_bus_aw_ready;
  wire                plicCtrl_io_bus_w_ready;
  wire                plicCtrl_io_bus_b_valid;
  wire       [1:0]    plicCtrl_io_bus_b_payload_resp;
  wire                plicCtrl_io_bus_ar_ready;
  wire                plicCtrl_io_bus_r_valid;
  wire       [31:0]   plicCtrl_io_bus_r_payload_data;
  wire       [1:0]    plicCtrl_io_bus_r_payload_resp;
  wire       [1:0]    plicCtrl_io_targets;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_payload;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_payload;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_payload;
  wire                integer_RfAllocationPlugin_logic_allocator_io_pop_ready;
  wire       [5:0]    integer_RfAllocationPlugin_logic_allocator_io_pop_values_0;
  wire                DataCachePlugin_logic_cache_io_load_cmd_ready;
  wire                DataCachePlugin_logic_cache_io_load_rsp_valid;
  wire       [31:0]   DataCachePlugin_logic_cache_io_load_rsp_payload_data;
  wire                DataCachePlugin_logic_cache_io_load_rsp_payload_fault;
  wire                DataCachePlugin_logic_cache_io_load_rsp_payload_redo;
  wire       [1:0]    DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlot;
  wire                DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlotAny;
  wire                DataCachePlugin_logic_cache_io_store_cmd_ready;
  wire                DataCachePlugin_logic_cache_io_store_rsp_valid;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_fault;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_redo;
  wire       [1:0]    DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlot;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlotAny;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_generationKo;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_flush;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_prefetch;
  wire       [31:0]   DataCachePlugin_logic_cache_io_store_rsp_payload_address;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_io;
  wire                DataCachePlugin_logic_cache_io_mem_read_cmd_valid;
  wire       [0:0]    DataCachePlugin_logic_cache_io_mem_read_cmd_payload_id;
  wire       [31:0]   DataCachePlugin_logic_cache_io_mem_read_cmd_payload_address;
  wire                DataCachePlugin_logic_cache_io_mem_read_rsp_ready;
  wire                DataCachePlugin_logic_cache_io_mem_write_cmd_valid;
  wire                DataCachePlugin_logic_cache_io_mem_write_cmd_payload_last;
  wire       [31:0]   DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_address;
  wire       [31:0]   DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_data;
  wire       [0:0]    DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_id;
  wire       [1:0]    DataCachePlugin_logic_cache_io_refillCompletions;
  wire                DataCachePlugin_logic_cache_io_refillEvent;
  wire                DataCachePlugin_logic_cache_io_writebackEvent;
  wire                DataCachePlugin_logic_cache_io_writebackBusy;
  wire                DataCachePlugin_logic_cache_io_tagEvent;
  wire                CommitPlugin_logic_free_lineEventStream_fifo_io_push_ready;
  wire                CommitPlugin_logic_free_lineEventStream_fifo_io_pop_valid;
  wire       [3:0]    CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_robId;
  wire       [0:0]    CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_mask;
  wire       [4:0]    CommitPlugin_logic_free_lineEventStream_fifo_io_occupancy;
  wire       [4:0]    CommitPlugin_logic_free_lineEventStream_fifo_io_availability;
  wire                EU0_DivPlugin_logic_div_io_cmd_ready;
  wire                EU0_DivPlugin_logic_div_io_rsp_valid;
  wire       [34:0]   EU0_DivPlugin_logic_div_io_rsp_payload_result;
  wire       [32:0]   EU0_DivPlugin_logic_div_io_rsp_payload_remain;
  wire                Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_valid;
  wire       [31:0]   Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_payload;
  wire                DispatchPlugin_logic_queue_io_push_ready;
  wire                DispatchPlugin_logic_queue_io_schedules_0_valid;
  wire       [7:0]    DispatchPlugin_logic_queue_io_schedules_0_payload_event;
  wire                DispatchPlugin_logic_queue_io_schedules_1_valid;
  wire       [7:0]    DispatchPlugin_logic_queue_io_schedules_1_payload_event;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_0_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_0_physRd;
  wire       [3:0]    DispatchPlugin_logic_queue_io_contexts_0_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_0_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_0_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_1_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_1_physRd;
  wire       [3:0]    DispatchPlugin_logic_queue_io_contexts_1_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_1_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_1_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_2_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_2_physRd;
  wire       [3:0]    DispatchPlugin_logic_queue_io_contexts_2_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_2_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_2_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_3_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_3_physRd;
  wire       [3:0]    DispatchPlugin_logic_queue_io_contexts_3_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_3_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_3_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_4_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_4_physRd;
  wire       [3:0]    DispatchPlugin_logic_queue_io_contexts_4_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_4_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_4_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_5_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_5_physRd;
  wire       [3:0]    DispatchPlugin_logic_queue_io_contexts_5_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_5_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_5_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_6_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_6_physRd;
  wire       [3:0]    DispatchPlugin_logic_queue_io_contexts_6_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_6_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_6_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_7_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_7_physRd;
  wire       [3:0]    DispatchPlugin_logic_queue_io_contexts_7_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_7_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_7_euCtx_1;
  wire       [7:0]    DispatchPlugin_logic_queue_io_usage;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_latches_io_reads_0_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_latches_io_reads_1_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_latches_io_reads_2_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_latches_io_reads_3_data;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_enable;
  wire       [3:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_rob;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_enable;
  wire       [3:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_rob;
  wire       [31:0]   _zz__zz_FetchPlugin_stages_1_MMU_IO;
  wire       [11:0]   _zz_FetchPlugin_stages_1_FETCH_ID;
  wire       [0:0]    _zz_FetchPlugin_stages_1_FETCH_ID_1;
  wire       [25:0]   _zz_FetchCachePlugin_logic_ways_0_mem_port;
  wire                _zz_FetchCachePlugin_logic_ways_0_mem_port_1;
  wire       [23:0]   _zz_FetchCachePlugin_logic_read_onWays_0_hits_bypassHits;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_usable;
  reg        [31:0]   _zz_AlignerPlugin_logic_extractors_0_pcWord;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_pcWord_1;
  wire       [29:0]   _zz_FrontendPlugin_aligned_PC_0;
  wire       [32:0]   _zz_BranchContextPlugin_logic_mem_earlyBranch_port;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push_1;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push_2;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push_3;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push_4;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_1;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_2;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_3;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_4;
  wire       [31:0]   _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port;
  wire       [48:0]   _zz_BtbPlugin_logic_mem_port;
  wire       [29:0]   _zz_BtbPlugin_logic_onLearn_port_payload_address;
  wire       [29:0]   _zz_BtbPlugin_logic_readCmd_entryAddress;
  wire       [1:0]    _zz_GSharePlugin_logic_mem_counter_port;
  wire       [6:0]    _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_1;
  wire       [23:0]   _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_2;
  wire       [6:0]    _zz_GSharePlugin_logic_onLearn_hash_1;
  wire       [23:0]   _zz_GSharePlugin_logic_onLearn_hash_2;
  wire       [4:0]    _zz_CommitPlugin_logic_ptr_allocNext;
  wire       [0:0]    _zz_CommitPlugin_logic_ptr_allocNext_1;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_commit_rowHit;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_age;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_0_age;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_1_age;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_2_age;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_3_age;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_4_age;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_1;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_2;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_3;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_4;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_5;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_6;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_7;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_8;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_9;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_10;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_11;
  wire       [0:0]    _zz_CommitPlugin_logic_reschedule_trap_5;
  wire       [0:0]    _zz_CommitPlugin_logic_reschedule_skipCommit;
  wire       [0:0]    _zz_CommitPlugin_logic_commit_active_1;
  wire       [0:0]    _zz_CommitPlugin_logic_commit_active_2;
  wire       [4:0]    _zz_CommitPlugin_logic_commit_head;
  wire       [3:0]    _zz_CommitPlugin_logic_free_robHit;
  wire       [31:0]   _zz_commit_pc_0_1;
  wire       [31:0]   _zz_commit_pc_0_2;
  reg        [0:0]    _zz_CommitDebugFilterPlugin_logic_commits;
  wire       [0:0]    _zz_CommitDebugFilterPlugin_logic_commits_1;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_0_value;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_0_value_1;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_0_value_2;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_0_value_3;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_1_value;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_1_value_1;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_1_value_2;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_1_value_3;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_2_value;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_2_value_1;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_2_value_2;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_2_value_3;
  wire       [31:0]   _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_1;
  wire       [31:0]   _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_2;
  wire       [11:0]   _zz__zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3;
  wire       [31:0]   _zz_ALU0_IntAluPlugin_logic_process_result;
  wire       [0:0]    _zz_ALU0_IntAluPlugin_logic_process_result_1;
  wire       [4:0]    _zz_ALU0_ShiftPlugin_logic_process_amplitude;
  wire       [31:0]   _zz_ALU0_ShiftPlugin_logic_process_reversed;
  wire                _zz_ALU0_ShiftPlugin_logic_process_reversed_1;
  wire       [0:0]    _zz_ALU0_ShiftPlugin_logic_process_reversed_2;
  wire       [20:0]   _zz_ALU0_ShiftPlugin_logic_process_reversed_3;
  wire                _zz_ALU0_ShiftPlugin_logic_process_reversed_4;
  wire       [0:0]    _zz_ALU0_ShiftPlugin_logic_process_reversed_5;
  wire       [9:0]    _zz_ALU0_ShiftPlugin_logic_process_reversed_6;
  wire       [32:0]   _zz_ALU0_ShiftPlugin_logic_process_shifted;
  wire       [32:0]   _zz_ALU0_ShiftPlugin_logic_process_shifted_1;
  wire       [31:0]   _zz_ALU0_ShiftPlugin_logic_process_patched;
  wire                _zz_ALU0_ShiftPlugin_logic_process_patched_1;
  wire       [0:0]    _zz_ALU0_ShiftPlugin_logic_process_patched_2;
  wire       [20:0]   _zz_ALU0_ShiftPlugin_logic_process_patched_3;
  wire                _zz_ALU0_ShiftPlugin_logic_process_patched_4;
  wire       [0:0]    _zz_ALU0_ShiftPlugin_logic_process_patched_5;
  wire       [9:0]    _zz_ALU0_ShiftPlugin_logic_process_patched_6;
  wire       [11:0]   _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [11:0]   _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_1;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4_1;
  wire       [29:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6_1;
  wire       [28:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8_1;
  wire       [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10_1;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12_1;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14_1;
  wire       [24:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16_1;
  wire       [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18_1;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20_1;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22_1;
  wire       [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24_1;
  wire       [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26_1;
  wire       [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28_1;
  wire       [17:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30_1;
  wire       [16:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32_1;
  wire       [15:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34_1;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36_1;
  wire       [13:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38_1;
  wire       [12:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40_1;
  wire       [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42_1;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44_1;
  wire       [9:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46_1;
  wire       [8:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48_1;
  wire       [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50_1;
  wire       [6:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52_1;
  wire       [5:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54_1;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56_1;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58_1;
  wire       [2:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60_1;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_63;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64;
  wire       [33:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_1;
  wire       [32:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_3;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_4;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_5;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_6;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_7;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_8;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_9;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_4;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_5;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_6;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_7;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_8;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_9;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_4;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_5;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_6;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_7;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_8;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_9;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_4;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_5;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_6;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_7;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_8;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_9;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_4;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_5;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_6;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_7;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_8;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_9;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_4;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_5;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_6;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_7;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_8;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_9;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_4;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_5;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_6;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_7;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_8;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_9;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_4;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_5;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_6;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_7;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_8;
  wire       [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_9;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_4;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_5;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_6;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_7;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_8;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_9;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_8;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_9;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_10;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_11;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_12;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_13;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_14;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_15;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_16;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_17;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_18;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_19;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_20;
  wire       [30:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_21;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_8;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_9;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_10;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_11;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_12;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_13;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_14;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_15;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_16;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_17;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_18;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_19;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_20;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_21;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_8;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_9;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_10;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_11;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_12;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_13;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_14;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_15;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_16;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_17;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_18;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_19;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_20;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_21;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_8;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_9;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_10;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_11;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_12;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_13;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_14;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_15;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_16;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_17;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_18;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_19;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_20;
  wire       [26:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_21;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_8;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_9;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_10;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_11;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_12;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_13;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_14;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_15;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_16;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_17;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_18;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_19;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_20;
  wire       [25:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_21;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_8;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_9;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_10;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_11;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_12;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_13;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_14;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_15;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_16;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_17;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_18;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_19;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_20;
  wire       [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_21;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_8;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_9;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_10;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_11;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_12;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_13;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_14;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_15;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_16;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_17;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_18;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_19;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_20;
  wire       [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_21;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_8;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_9;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_10;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_11;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_12;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_13;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_14;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_15;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_16;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_17;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_18;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_19;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_20;
  wire       [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_21;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_7;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_8;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_9;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_10;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_11;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_12;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_13;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_14;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_15;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_16;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_17;
  wire       [69:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_18;
  wire       [34:0]   _zz_EU0_DivPlugin_logic_rsp_selected;
  wire       [34:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_1;
  wire       [34:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_2;
  wire       [34:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_3;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_4;
  wire       [20:0]   _zz_EU0_BranchPlugin_logic_process_target_b;
  wire       [11:0]   _zz_EU0_BranchPlugin_logic_process_target_b_1;
  wire       [12:0]   _zz_EU0_BranchPlugin_logic_process_target_b_2;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
  wire       [1:0]    _zz_EU0_BranchPlugin_logic_process_slices;
  wire       [0:0]    _zz_EU0_BranchPlugin_logic_process_slices_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1;
  wire       [31:0]   _zz_LsuPlugin_peripheralBus_toAxiLite4_addr;
  wire       [2:0]    _zz_BranchContextPlugin_logic_onCommit_commitedNext;
  reg        [0:0]    _zz_BranchContextPlugin_logic_onCommit_commitedNext_1;
  wire       [0:0]    _zz_BranchContextPlugin_logic_onCommit_commitedNext_2;
  wire       [24:0]   _zz_HistoryPlugin_logic_onCommit_valueNext_1;
  wire       [24:0]   _zz_HistoryPlugin_logic_update_pushes_0_stateNext_1;
  wire       [24:0]   _zz_HistoryPlugin_logic_update_pushes_2_stateNext_1;
  wire       [23:0]   _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_1;
  wire       [23:0]   _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_2;
  wire       [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_1;
  wire       [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_2;
  wire       [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_1;
  wire       [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_2;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_healPush_1;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_healPush_2;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_tracker_freeNext;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_tracker_freeNext_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_tracker_freeNext_2;
  reg        [0:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount_1;
  wire       [2:0]    _zz_when_Lsu2Plugin_l454;
  wire       [2:0]    _zz_when_Lsu2Plugin_l454_1;
  wire       [2:0]    _zz_when_Lsu2Plugin_l454_2;
  wire       [2:0]    _zz_when_Lsu2Plugin_l454_3;
  wire       [2:0]    _zz_when_Lsu2Plugin_l454_4;
  wire       [2:0]    _zz_when_Lsu2Plugin_l454_5;
  wire       [2:0]    _zz_when_Lsu2Plugin_l454_6;
  wire       [2:0]    _zz_when_Lsu2Plugin_l454_7;
  wire       [6:0]    _zz_Lsu2Plugin_logic_lq_onCommit_priority_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_onCommit_free_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_onCommit_free_1_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_ptr_free;
  wire       [21:0]   _zz_Lsu2Plugin_logic_lq_hazardPrediction_mem_port;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_hitPrediction_mem_port;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext_2;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext_3;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext_4;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1_1;
  reg        [0:0]    _zz_Lsu2Plugin_logic_allocation_loads_requestsCount;
  wire       [0:0]    _zz_Lsu2Plugin_logic_allocation_loads_requestsCount_1;
  reg        [0:0]    _zz_Lsu2Plugin_logic_allocation_stores_requestsCount;
  wire       [0:0]    _zz_Lsu2Plugin_logic_allocation_stores_requestsCount_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_sqAlloc_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_doSpecial_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_doSpecial_port;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_lqAlloc_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_feededOnce_port;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_addressPre_port;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_addressPre_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_physRd_port;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_physRd_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_robId_port;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_robId_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_pc_port;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_pc_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_writeRd_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_writeRd_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_lr_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_lr_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_size_port;
  wire       [1:0]    _zz_Lsu2Plugin_logic_lq_mem_size_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_unsigned_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_unsigned_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_needTranslation_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_needTranslation_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_addressPre_port;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPre_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_robId_port;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_robId_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_amo_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_amo_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_sc_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_sc_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_size_port;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sq_mem_size_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_needTranslation_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_needTranslation_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_data_port;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port_1;
  wire       [7:0]    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh;
  wire       [7:0]    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lqSqArbitration_s1_cmp;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_sqAlloc_port_1;
  wire       [3:0]    _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT;
  wire       [3:0]    _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_feededOnce_port_1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_3;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_3;
  wire       [7:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_addressPost_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_io_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_needTranslation_port_2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPost_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_io_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_needTranslation_port_2;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_3;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_3;
  wire       [7:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh;
  reg        [7:0]    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_1;
  reg        [7:0]    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_3;
  reg                 _zz__zz_when_Lsu2Plugin_l1348;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_doSpecial_port_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_doSpecial_port_1;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_1;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_2;
  wire       [1:0]    _zz_when_SInt_l132;
  wire       [0:0]    _zz_when_SInt_l138;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_ptr_writeBack;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_ptr_writeBack_1;
  wire       [2:0]    _zz_Lsu2Plugin_setup_specialTrap_payload_cause;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_3;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_4;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_5;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_6;
  wire       [1:0]    _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_7;
  wire       [31:0]   _zz_EU0_BranchPlugin_setup_intFormatPort_payload;
  wire       [4:0]    _zz_EU0_BranchPlugin_setup_reschedule_payload_reason;
  wire       [64:0]   _zz_BranchContextPlugin_logic_mem_finalBranch_port;
  wire       [31:0]   _zz_EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice;
  wire       [1:0]    _zz_EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1;
  wire       [44:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port_1;
  wire       [44:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port_1;
  wire       [44:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port_1;
  wire       [44:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port_1;
  wire       [1:0]    _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
  wire       [0:0]    _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1;
  wire       [24:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port_1;
  wire       [24:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port_1;
  wire       [44:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port_1;
  wire       [44:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port_1;
  wire       [44:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port_1;
  wire       [44:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port_1;
  wire       [1:0]    _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
  wire       [0:0]    _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1;
  wire       [24:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port_1;
  wire       [24:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_6;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_1;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_3;
  wire       [11:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_4;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_5;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_6;
  wire       [11:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_7;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_8;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_9;
  wire       [11:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_10;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_11;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_12;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_13;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault;
  wire       [2:0]    _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  reg        [2:0]    _zz_CsrRamPlugin_logic_writeLogic_port_payload_address;
  reg        [31:0]   _zz_CsrRamPlugin_logic_writeLogic_port_payload_data;
  wire       [1:0]    _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  reg        [2:0]    _zz_CsrRamPlugin_logic_readLogic_port_address;
  wire       [0:0]    _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented;
  wire       [12:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_1;
  wire       [0:0]    _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_2;
  wire       [1:0]    _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_3;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_setup_onDecodeAddress;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_setup_onReadAddress;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [4:0]    _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_setup_onWriteAddress;
  wire       [31:0]   _zz_csrAccess_payload_address;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_6;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineException;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_1;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_2;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_3;
  wire       [11:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_4;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_5;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_6;
  wire       [11:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_7;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_8;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_9;
  wire       [11:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_10;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_11;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_12;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_13;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault;
  wire       [1:0]    _zz_MmuPlugin_logic_refill_portsRequests_ohFirst_masked;
  wire       [3:0]    _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask_1;
  wire       [3:0]    _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask_1;
  wire       [1:0]    _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask;
  wire       [1:0]    _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_2;
  wire                _zz_FrontendPlugin_decoded_LEGAL_0_3;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_4;
  wire       [18:0]   _zz_FrontendPlugin_decoded_LEGAL_0_5;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_6;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_7;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_8;
  wire                _zz_FrontendPlugin_decoded_LEGAL_0_9;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_10;
  wire       [12:0]   _zz_FrontendPlugin_decoded_LEGAL_0_11;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_12;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_13;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_14;
  wire                _zz_FrontendPlugin_decoded_LEGAL_0_15;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_16;
  wire       [6:0]    _zz_FrontendPlugin_decoded_LEGAL_0_17;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_18;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_19;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_20;
  wire                _zz_FrontendPlugin_decoded_LEGAL_0_21;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_22;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_23;
  wire       [0:0]    _zz_FrontendPlugin_decoded_READ_RS_0_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_READ_RS_1_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_WRITE_RD_0_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_0_2;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_0_3;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_0_4;
  wire                _zz_FrontendPlugin_decoded_WRITE_RD_0_5;
  wire                _zz_FrontendPlugin_decoded_WRITE_RD_0_6;
  wire       [0:0]    _zz_FrontendPlugin_decoded_ALU0_SEL_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_EU0_SEL_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LQ_ALLOC_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_SQ_ALLOC_0_2;
  wire       [0:0]    _zz_DecoderPlugin_logic_exception_compressedFault;
  wire       [0:0]    _zz_DecoderPlugin_logic_exception_fetchFault;
  wire       [0:0]    _zz_DecoderPlugin_logic_exception_fetchFaultPage;
  wire       [0:0]    _zz_DecoderPlugin_logic_exception_debugEnter;
  wire       [31:0]   _zz_DecoderPlugin_setup_exceptionPort_payload_tval;
  wire       [31:0]   _zz_DecoderPlugin_setup_exceptionPort_payload_tval_1;
  wire       [1:0]    _zz_DecoderPlugin_setup_exceptionPort_payload_tval_2;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_4;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_5;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0_1;
  wire       [11:0]   _zz_FrontendPlugin_decoded_OP_ID;
  wire       [0:0]    _zz_FrontendPlugin_decoded_OP_ID_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_JAL_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_JALR_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_ANY_0;
  wire       [12:0]   _zz__zz_FrontendPlugin_decoded_OFFSET_0;
  wire       [20:0]   _zz__zz_FrontendPlugin_decoded_OFFSET_0_1;
  wire       [1:0]    _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_INC_0;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_INC_0_1;
  wire       [3:0]    _zz_FrontendPlugin_decoded_PC_INC_0_2;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2;
  wire       [5:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1;
  wire       [5:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2;
  wire       [5:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1;
  wire       [5:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_1;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_2;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_2;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_1;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_2;
  wire       [1:0]    _zz_BranchContextPlugin_free_learn_GSHARE_COUNTER_0;
  wire       [3:0]    _zz_DispatchPlugin_logic_ptr_next;
  wire       [7:0]    _zz_DispatchPlugin_logic_push_slots_0_events_0;
  wire       [2:0]    _zz_DispatchPlugin_logic_push_slots_0_events_0_1;
  wire       [3:0]    _zz_DispatchPlugin_logic_push_slots_0_events_0_2;
  wire       [7:0]    _zz_DispatchPlugin_logic_push_slots_0_events_1;
  wire       [2:0]    _zz_DispatchPlugin_logic_push_slots_0_events_1_1;
  wire       [3:0]    _zz_DispatchPlugin_logic_push_slots_0_events_1_2;
  wire       [3:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID;
  wire       [3:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID;
  wire       [3:0]    _zz_DispatchPlugin_logic_wake_dynamic_offseted_0_payload;
  wire       [3:0]    _zz_DispatchPlugin_logic_wake_dynamic_offseted_1_payload;
  wire       [3:0]    _zz_DispatchPlugin_logic_wake_dynamic_offseted_2_payload;
  wire       [3:0]    _zz_DispatchPlugin_logic_wake_dynamic_offseted_3_payload;
  wire       [7:0]    _zz_DispatchPlugin_logic_wake_dynamic_masks_0;
  wire       [7:0]    _zz_DispatchPlugin_logic_wake_dynamic_masks_1;
  wire       [7:0]    _zz_DispatchPlugin_logic_wake_dynamic_masks_2;
  wire       [7:0]    _zz_DispatchPlugin_logic_wake_dynamic_masks_3;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_0_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_1_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_2_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_3_port;
  wire       [0:0]    _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_1;
  wire       [0:0]    _zz_integer_RfAllocationPlugin_logic_push_mask_0_1;
  wire       [0:0]    _zz_integer_RfAllocationPlugin_logic_push_mask_0_2;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_PC_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port_1;
  wire       [0:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1;
  wire       [0:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_2;
  wire       [0:0]    _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1;
  wire       [0:0]    _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_2;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_1;
  wire       [5:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_1;
  wire       [5:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2;
  wire       [5:0]    _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_1;
  wire       [5:0]    _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2;
  wire       [4:0]    _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_1;
  wire       [4:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_1;
  wire       [4:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_1;
  wire       [5:0]    _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_1;
  wire       [5:0]    _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_1;
  wire       [0:0]    _zz_BranchContextPlugin_logic_onCommit_isBranch_0_1;
  wire       [0:0]    _zz_BranchContextPlugin_logic_onCommit_isBranch_0_2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port_1;
  wire       [0:0]    _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1;
  wire       [0:0]    _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_port_1;
  wire       [0:0]    _zz_HistoryPlugin_logic_onCommit_isTaken_0_1;
  wire       [0:0]    _zz_HistoryPlugin_logic_onCommit_isTaken_0_2;
  wire                _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port;
  wire       [3:0]    _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2;
  wire                _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port_1;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port_1;
  wire       [1:0]    _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port_1;
  wire       [3:0]    _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port_1;
  wire       [6:0]    _zz_PcPlugin_logic_init_counter;
  wire       [0:0]    _zz_PcPlugin_logic_init_counter_1;
  wire       [31:0]   _zz_PcPlugin_logic_fetchPc_pc;
  wire       [2:0]    _zz_PcPlugin_logic_fetchPc_pc_1;
  wire       [31:0]   _zz_PrivilegedPlugin_setup_ramWrite_data;
  wire       [31:0]   _zz_PrivilegedPlugin_setup_ramWrite_data_1;
  wire       [31:0]   _zz_PrivilegedPlugin_logic_readed;
  wire       [31:0]   _zz_PrivilegedPlugin_logic_readed_1;
  wire       [3:0]    _zz_PrivilegedPlugin_logic_readed_2;
  wire       [3:0]    _zz_PrivilegedPlugin_logic_readed_3;
  wire       [1:0]    _zz_PrivilegedPlugin_logic_readed_4;
  wire       [1:0]    _zz_PrivilegedPlugin_logic_readed_5;
  wire       [0:0]    _zz_PrivilegedPlugin_logic_readed_6;
  wire                FetchPlugin_stages_2_isFlushingRoot;
  wire                FetchPlugin_stages_1_isFlushingRoot;
  wire                FetchPlugin_stages_0_isFlushed;
  wire                FetchPlugin_stages_1_isFlushingNext;
  wire                FetchPlugin_stages_1_isThrown;
  wire                FetchPlugin_stages_2_isFlushed;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_FETCH_PC_INC;
  reg        [1:0]    FetchPlugin_stages_2_GSHARE_COUNTER_0;
  reg                 FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE;
  reg                 FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID;
  reg        [31:0]   FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT;
  reg        [0:0]    FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT;
  reg                 FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID;
  reg        [23:0]   FetchPlugin_stages_1_BRANCH_HISTORY;
  reg        [11:0]   FetchPlugin_stages_2_FETCH_ID;
  reg        [31:0]   FetchPlugin_stages_1_Fetch_FETCH_PC_INC;
  wire                FrontendPlugin_dispatch_isFlushingRoot;
  wire                FrontendPlugin_decoded_isFlushingRoot;
  wire                FrontendPlugin_decompressed_isFlushed;
  wire                FrontendPlugin_allocated_isFlushed;
  wire                FrontendPlugin_dispatch_isFlushed;
  wire                FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_0;
  wire                FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_0;
  wire                FrontendPlugin_allocated_EU0_SEL_0;
  reg                 FrontendPlugin_serialized_EU0_SEL_0;
  wire                FrontendPlugin_allocated_ALU0_SEL_0;
  reg                 FrontendPlugin_serialized_ALU0_SEL_0;
  wire                FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_0;
  wire                FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_0;
  wire       [1:0]    FrontendPlugin_allocated_GSHARE_COUNTER_0_0;
  reg        [1:0]    FrontendPlugin_serialized_GSHARE_COUNTER_0_0;
  wire       [1:0]    FrontendPlugin_decoded_GSHARE_COUNTER_0_0;
  wire                FrontendPlugin_allocated_Prediction_IS_BRANCH_0;
  wire                FrontendPlugin_allocated_SQ_ALLOC_0;
  reg                 FrontendPlugin_serialized_SQ_ALLOC_0;
  wire                FrontendPlugin_allocated_LQ_ALLOC_0;
  reg                 FrontendPlugin_serialized_LQ_ALLOC_0;
  reg        [11:0]   FrontendPlugin_serialized_OP_ID;
  reg        [23:0]   FrontendPlugin_serialized_BRANCH_HISTORY_0;
  wire       [23:0]   FrontendPlugin_decoded_BRANCH_HISTORY_0;
  wire       [23:0]   FrontendPlugin_decompressed_BRANCH_HISTORY_0;
  reg                 FrontendPlugin_serialized_READ_RS_1_0;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RS_1_0;
  reg                 FrontendPlugin_serialized_READ_RS_0_0;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RS_0_0;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RD_0;
  reg        [31:0]   FrontendPlugin_serialized_PC_0;
  reg                 FrontendPlugin_serialized_WRITE_RD_0;
  reg        [11:0]   FrontendPlugin_serialized_FETCH_ID_0;
  wire                FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_0;
  wire                FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_0;
  wire       [31:0]   FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  wire       [31:0]   FrontendPlugin_decompressed_PC_0;
  wire                FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_0;
  wire                FrontendPlugin_decompressed_Frontend_FETCH_FAULT_0;
  wire                FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_0;
  wire       [11:0]   FrontendPlugin_decompressed_FETCH_ID_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0;
  reg                 FrontendPlugin_dispatch_READ_RS_1_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0;
  reg                 FrontendPlugin_dispatch_READ_RS_0_0;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 _zz_3;
  reg                 _zz_4;
  reg                 _zz_5;
  wire                DispatchPlugin_logic_pop_1_stagesList_0_isFlushed;
  wire                DispatchPlugin_logic_pop_1_stagesList_1_isFlushed;
  reg                 DispatchPlugin_logic_pop_1_stagesList_1_ready;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_0;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_1;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_2;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_3;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RS_1;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_0;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_1;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_2;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_3;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_0;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_1;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_2;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_3;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RS_0;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_0;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_1;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_2;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_3;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_0;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_1;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_2;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_3;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RD;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_0;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_1;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_2;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_3;
  wire                DispatchPlugin_logic_pop_1_stagesList_0_LATENCY_0;
  reg        [3:0]    DispatchPlugin_logic_pop_1_stagesList_1_OFFSET;
  reg        [2:0]    DispatchPlugin_logic_pop_1_stagesList_1_UINT;
  wire       [3:0]    DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID;
  wire       [2:0]    DispatchPlugin_logic_pop_1_stagesList_0_UINT;
  wire                DispatchPlugin_logic_pop_1_stagesList_0_ready;
  wire       [3:0]    DispatchPlugin_logic_pop_1_stagesList_0_OFFSET;
  wire       [7:0]    DispatchPlugin_logic_pop_1_stagesList_0_OH;
  wire                DispatchPlugin_logic_pop_0_stagesList_0_isFlushed;
  wire                DispatchPlugin_logic_pop_0_stagesList_1_isFlushed;
  reg                 DispatchPlugin_logic_pop_0_stagesList_1_LATENCY_0;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_0;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_1;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_2;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_3;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_PHYS_RD;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3;
  wire                DispatchPlugin_logic_pop_0_stagesList_0_LATENCY_0;
  reg        [3:0]    DispatchPlugin_logic_pop_0_stagesList_1_OFFSET;
  reg        [2:0]    DispatchPlugin_logic_pop_0_stagesList_1_UINT;
  wire       [3:0]    DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID;
  wire       [2:0]    DispatchPlugin_logic_pop_0_stagesList_0_UINT;
  wire                DispatchPlugin_logic_pop_0_stagesList_0_ready;
  wire       [3:0]    DispatchPlugin_logic_pop_0_stagesList_0_OFFSET;
  wire       [7:0]    DispatchPlugin_logic_pop_0_stagesList_0_OH;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RS_1_0;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RS_0_0;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RD_0;
  reg                 FrontendPlugin_dispatch_EU0_SEL_0;
  reg                 FrontendPlugin_dispatch_ALU0_SEL_0;
  wire                FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_0;
  wire       [3:0]    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0;
  wire                FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_0;
  wire       [3:0]    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0;
  reg                 FrontendPlugin_dispatch_WRITE_RD_0;
  reg                 FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_0;
  reg                 FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_0;
  reg        [1:0]    FrontendPlugin_dispatch_GSHARE_COUNTER_0_0;
  reg        [23:0]   FrontendPlugin_dispatch_BRANCH_HISTORY_0;
  reg        [1:0]    FrontendPlugin_dispatch_BRANCH_ID_0;
  reg                 FrontendPlugin_dispatch_BRANCH_SEL_0;
  reg                 _zz_6;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_isFlushed;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_1_isFlushed;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_isThrown;
  wire                EU0_ExecutionUnitBase_pipeline_execute_1_isFlushed;
  wire                EU0_ExecutionUnitBase_pipeline_execute_2_isFlushed;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E2;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E2;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E2;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_execute_1_PHYS_RD;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_WRITE_RD;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_Frontend_MICRO_OP;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_PC_FALSE;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_CsrAccessPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_WFI;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_WFI;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_WFI;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_VMA;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_VMA;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_VMA;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FLUSH_DATA;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FLUSH_DATA;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FLUSH_DATA;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_I;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_I;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_I;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_XRET;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_XRET;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_XRET;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_ECALL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_ECALL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_ECALL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_EBREAK;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_EBREAK;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_EBREAK;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_HIGH;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_HIGH;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_HIGH;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_CLEAR;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_MASK;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_IMM;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LOAD;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LR;
  reg        [3:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_LSU_ID;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_AMO;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SC;
  reg        [0:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_MSB;
  reg        [3:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SEL;
  reg        [1:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_PC;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP;
  reg        [1:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_REM;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS2_SIGNED;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS1_SIGNED;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS2;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS1;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_completion_SEL_E2;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_execute_2_PHYS_RD;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL;
  wire       [1:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL;
  wire       [0:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID;
  wire       [1:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_ready;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_isFlushed;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_1_isFlushed;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_isFlushed;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0;
  reg        [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  reg        [3:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL;
  reg        [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL;
  reg        [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_ready;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  wire       [3:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
  wire       [3:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  reg                 FrontendPlugin_dispatch_Prediction_IS_BRANCH_0;
  reg                 FrontendPlugin_serialized_Prediction_IS_BRANCH_0;
  wire                FrontendPlugin_serialized_isFlushed;
  wire                FrontendPlugin_serialized_ready;
  wire       [3:0]    FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_0;
  reg                 FrontendPlugin_serialized_RAS_POP_0;
  reg                 DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_1;
  reg                 FrontendPlugin_serialized_RAS_PUSH_0;
  wire                FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0;
  reg        [31:0]   FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  reg                 FrontendPlugin_serialized_BRANCH_EARLY_0_taken;
  reg        [31:0]   FrontendPlugin_serialized_BRANCH_EARLY_0_pc;
  wire                FrontendPlugin_serialized_BRANCH_SEL_0;
  reg                 FrontendPlugin_serialized_CAN_IMPROVE_0;
  reg                 FrontendPlugin_serialized_Frontend_DECODED_MASK_0;
  wire                FrontendPlugin_serialized_NEED_CORRECTION_0;
  wire                FrontendPlugin_serialized_MISSMATCH_0;
  wire                FrontendPlugin_serialized_MISSMATCH_HISTORY_0;
  reg                 FrontendPlugin_serialized_BAD_RET_PC_0;
  wire                FrontendPlugin_serialized_MISSMATCH_PC_0;
  reg                 FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0;
  reg                 FrontendPlugin_serialized_IS_ANY_0;
  reg        [31:0]   FrontendPlugin_serialized_PC_INC_0;
  reg                 FrontendPlugin_serialized_BRANCHED_PREDICTION_0;
  wire       [31:0]   FrontendPlugin_serialized_PC_PREDICTION_0;
  reg                 FrontendPlugin_serialized_IS_JALR_0;
  reg        [31:0]   FrontendPlugin_serialized_PC_TARGET_PRE_RAS_0;
  reg        [31:0]   FrontendPlugin_serialized_PC_TARGET_0;
  wire                FrontendPlugin_decoded_BRANCHED_PREDICTION_0;
  wire                FrontendPlugin_decoded_CAN_IMPROVE_0;
  wire       [31:0]   FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  wire                FrontendPlugin_decoded_BAD_RET_PC_0;
  wire       [31:0]   FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0;
  wire       [31:0]   FrontendPlugin_decoded_PC_INC_0;
  wire       [0:0]    FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_0;
  wire                FrontendPlugin_decoded_CONDITIONAL_PREDICTION_0;
  wire                FrontendPlugin_decoded_RAS_POP_0;
  wire                FrontendPlugin_decoded_RAS_PUSH_0;
  wire       [31:0]   FrontendPlugin_decoded_OFFSET_0;
  wire                FrontendPlugin_decoded_IS_ANY_0;
  wire                FrontendPlugin_decoded_Prediction_IS_BRANCH_0;
  wire                FrontendPlugin_decoded_IS_JALR_0;
  reg        [31:0]   FrontendPlugin_dispatch_Frontend_MICRO_OP_0;
  wire                FrontendPlugin_dispatch_LATENCY_0_0;
  wire       [11:0]   FrontendPlugin_allocated_OP_ID /* verilator public */ ;
  reg        [11:0]   FrontendPlugin_decoded_OP_ID /* verilator public */ ;
  wire       [3:0]    FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_0;
  wire       [31:0]   FrontendPlugin_allocated_Frontend_MICRO_OP_0;
  wire                FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0;
  wire                FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0;
  wire                FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0;
  wire                FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0;
  reg        [31:0]   FrontendPlugin_serialized_Frontend_MICRO_OP_0;
  wire                FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_0;
  wire       [31:0]   FrontendPlugin_decoded_PC_0 /* verilator public */ ;
  wire                FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_0;
  wire                FrontendPlugin_decoded_isFlushed;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RS_1_0;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RS_0_0;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RD_0;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_MICRO_OP_0;
  wire                FrontendPlugin_decoded_Frontend_DECODED_MASK_0 /* verilator public */ ;
  wire                FrontendPlugin_decoded_Frontend_FETCH_FAULT_0;
  wire                FrontendPlugin_decoded_Frontend_MASK_ALIGNED_0;
  wire                FrontendPlugin_decoded_TRAP_0;
  wire                FrontendPlugin_decoded_SQ_ALLOC_0;
  wire                FrontendPlugin_decoded_LQ_ALLOC_0;
  wire                FrontendPlugin_decoded_EU0_SEL_0;
  wire                FrontendPlugin_decoded_ALU0_SEL_0;
  wire                FrontendPlugin_decoded_WRITE_RD_0;
  wire                FrontendPlugin_decoded_READ_RS_1_0;
  wire                FrontendPlugin_decoded_READ_RS_0_0;
  wire                FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_0;
  wire                FrontendPlugin_decoded_LEGAL_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_isFlushed;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_isThrown;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_isFlushed;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_isThrown;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_isFlushed;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_isThrown;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_isFlushed;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_isFlushed;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_isFlushed;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH_PC;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH_PC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_SP_FP_ADDRESS;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_SP_FP_ADDRESS;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION_COUNTER;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION_COUNTER;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_AMO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_AMO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_SC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_SC;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_DELTA;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_DELTA;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_VALID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_VALID;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SCORE;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SCORE;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_MMU_TRANSLATED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LR;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LR;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_SQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_1_PHYS_RD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_WRITE_RD;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_ROB_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_UNSIGNED;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_1_SIZE;
  reg                 FetchPlugin_stages_1_MMU_ACCESS_FAULT;
  reg                 FetchPlugin_stages_1_MMU_PAGE_FAULT;
  reg                 FetchPlugin_stages_1_MMU_ALLOW_WRITE;
  reg                 FetchPlugin_stages_1_MMU_ALLOW_READ;
  reg                 FetchPlugin_stages_1_MMU_ALLOW_EXECUTE;
  reg                 FetchPlugin_stages_1_MMU_REDO;
  reg        [31:0]   FetchPlugin_stages_1_MMU_TRANSLATED;
  wire                FetchPlugin_stages_1_MMU_IO;
  reg        [1:0]    FetchPlugin_stages_1_MMU_L1_HITS;
  reg        [1:0]    FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_pageFault;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_accessFault;
  wire       [7:0]    FetchPlugin_stages_1_MMU_L1_ENTRIES_0_virtualAddress;
  wire       [9:0]    FetchPlugin_stages_1_MMU_L1_ENTRIES_0_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowRead;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowUser;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_pageFault;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_accessFault;
  wire       [7:0]    FetchPlugin_stages_1_MMU_L1_ENTRIES_1_virtualAddress;
  wire       [9:0]    FetchPlugin_stages_1_MMU_L1_ENTRIES_1_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowRead;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowUser;
  reg        [3:0]    FetchPlugin_stages_1_MMU_L0_HITS;
  reg        [3:0]    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_pageFault;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_accessFault;
  wire       [17:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_0_virtualAddress;
  wire       [19:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_0_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowRead;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowUser;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_pageFault;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_accessFault;
  wire       [17:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_1_virtualAddress;
  wire       [19:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_1_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowRead;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowUser;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_pageFault;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_accessFault;
  wire       [17:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_2_virtualAddress;
  wire       [19:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_2_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowRead;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowUser;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_pageFault;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_accessFault;
  wire       [17:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_3_virtualAddress;
  wire       [19:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_3_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowRead;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowUser;
  wire                FetchPlugin_stages_1_isRemoved;
  wire                FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded;
  wire                FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_0;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_1;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_2;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_3;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_4;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_5;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_OH;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_MMU_BYPASS_TRANSLATION;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_WRITE;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_EXECUTE;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_2_PC;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_2_Frontend_MICRO_OP;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_ready;
  reg        [3:0]    EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_CLEAR;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_IMM;
  reg                 _zz_7;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_accessFault;
  reg        [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_virtualAddress;
  reg        [9:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_accessFault;
  reg        [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_virtualAddress;
  reg        [9:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowUser;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS_PRE_VALID;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_HITS_PRE_VALID;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_accessFault;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_virtualAddress;
  wire       [9:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_accessFault;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_virtualAddress;
  wire       [9:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_accessFault;
  reg        [17:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_virtualAddress;
  reg        [19:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_accessFault;
  reg        [17:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_virtualAddress;
  reg        [19:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_accessFault;
  reg        [17:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_virtualAddress;
  reg        [19:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_accessFault;
  reg        [17:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_virtualAddress;
  reg        [19:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowUser;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_accessFault;
  wire       [17:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_virtualAddress;
  wire       [19:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_accessFault;
  wire       [17:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_virtualAddress;
  wire       [19:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_accessFault;
  wire       [17:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_virtualAddress;
  wire       [19:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_accessFault;
  wire       [17:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_virtualAddress;
  wire       [19:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_isRemoved;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_isRemoved;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL_overloaded;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_PC_TRUE;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_PC;
  reg        [1:0]    EU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID;
  reg                 _zz_8;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  reg        [1:0]    EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  reg        [3:0]    EU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET;
  wire                EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_pc;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_2_PC_FALSE;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET;
  reg                 _zz_FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH_PC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_SP_FP_ADDRESS;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION_COUNTER;
  reg                 _zz_9;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_AMO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_SC;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ROB;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_DELTA;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_VALID;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE;
  reg                 _zz_10;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_MMU_TRANSLATED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LR;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_WRITE_RD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_IS_IO;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_resulting;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_resulting;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_WAIT_FEED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_ready;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_CTRL;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_valid;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_data;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_fault;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlot;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlotAny;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_ADDRESS_PRE_TRANSLATION;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_3_PHYS_RD;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ID;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_valid;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_data;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_fault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_redo;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlot;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_valid;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_data;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_fault;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlot;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_valid;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_data;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_fault;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlot;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_TRAP_SPECULATION;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_CTRL;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_WRITE;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_PAGE_FAULT;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_MISS_ALIGNED;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_WRITE_FAILURE;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_2_PHYS_RD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_ACCESS_FAULT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_READ;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_WRITE_RD;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_LQ_ID;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_REDO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_IS_IO;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_ready;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_HIT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_UNSIGNED;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_valid;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_fault;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlot;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlotAny;
  wire       [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ID;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_RESCHEDULE;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ROB;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_NO_YOUNGER;
  reg        [7:0]    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER;
  reg        [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_BYPASS_SUCCESS;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_2_SIZE;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_TRANSLATED;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_overloaded;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED_overloaded;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED;
  reg                 _zz_11;
  reg                 _zz_12;
  reg                 _zz_13;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID;
  reg                 _zz_14;
  reg                 _zz_15;
  reg                 _zz_16;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_ready;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_OH;
  wire       [2:0]    Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_ID;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_HIT;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_NO_OLDER;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_TRANSLATED_AS_IO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_IS_IO;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_POST_TRANSLATION;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION;
  reg                 _zz_17;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH_PC;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SQID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SQID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SQID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_FEEDED;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT;
  wire       [2:0]    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SQID;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_feed_SQ_PTR_FREE;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_SQCHECK_END_ID;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_LQCHECK_START_ID;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD_agu;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD_agu;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_agu;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_SP_FP_ADDRESS;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION_COUNTER;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_SC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_AMO;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SCORE;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_LR;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_UNSIGNED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_store;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_load;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_store;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_load;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_0_SIZE;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_0_SIZE_store;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_0_SIZE_load;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_store;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_load;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_store;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_load;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s1_ready;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_isRemoved;
  reg                 _zz_Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_ready;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_stages_0_SQ_ROB_FULL;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_stages_0_LQ_ROB_FULL;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ;
  reg        [2:0]    Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID;
  reg        [2:0]    Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s1_LQ_HIT;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s1_SQ_HIT;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_LQ_OLDER_THAN_SQ;
  reg        [4:0]    Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ROB_FULL;
  reg        [4:0]    Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ROB_FULL;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_ready;
  wire       [4:0]    Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ROB_FULL;
  wire       [4:0]    Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ROB_FULL;
  wire       [2:0]    Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID;
  wire       [2:0]    Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH;
  reg        [3:0]    FrontendPlugin_dispatch_ROB_ID /* verilator public */ ;
  reg        [3:0]    Lsu2Plugin_logic_allocation_stores_alloc_1;
  reg                 _zz_18;
  reg                 _zz_19;
  reg                 _zz_20;
  reg        [3:0]    Lsu2Plugin_logic_allocation_loads_alloc_1;
  reg                 _zz_21;
  reg        [4:0]    FrontendPlugin_dispatch_ARCH_RS_0_0;
  reg                 _zz_22;
  reg                 _zz_23;
  reg                 FrontendPlugin_dispatch_ready;
  wire       [2:0]    FrontendPlugin_dispatch_SQ_ID_0;
  wire       [2:0]    FrontendPlugin_dispatch_LQ_ID_0;
  reg                 FrontendPlugin_dispatch_SQ_ALLOC_0;
  reg                 FrontendPlugin_dispatch_LQ_ALLOC_0;
  reg                 FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 /* verilator public */ ;
  reg        [3:0]    FrontendPlugin_dispatch_LSU_ID_0;
  reg        [3:0]    Lsu2Plugin_logic_sq_onCommit_commitComb_1;
  reg                 _zz_24;
  reg                 _zz_25;
  reg        [3:0]    Lsu2Plugin_logic_lq_onCommit_free_1;
  reg        [6:0]    Lsu2Plugin_logic_lq_onCommit_priority_1;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 /* verilator public */ ;
  wire                FrontendPlugin_decoded_IS_JAL_0;
  wire       [23:0]   FrontendPlugin_allocated_BRANCH_HISTORY_0 /* verilator public */ ;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_2_stateNext_1;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_0_stateNext_1;
  reg        [23:0]   HistoryPlugin_logic_onCommit_valueNext_1;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RS_1_0;
  wire                FrontendPlugin_allocated_READ_RS_1_0;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RS_1_0;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RS_0_0;
  wire                FrontendPlugin_allocated_READ_RS_0_0;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RS_0_0;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RD_FREE_0;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RD_0;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_WFI;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LOAD;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LR;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_execute_0_LSU_ID;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_AMO;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SC;
  wire       [0:0]    EU0_ExecutionUnitBase_pipeline_execute_0_ROB_MSB;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_isRemoved;
  wire       [1:0]    EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_PC_TARGET;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_PC;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
  wire       [1:0]    EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_BranchPlugin_SEL;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_DIV_RESULT;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_DIV_REVERT_RESULT;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_REM;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_ready;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_0_ready;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_DIV_REVERT_RESULT;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_HIGH;
  wire       [69:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0;
  reg        [2:0]    EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_7;
  reg        [14:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_6;
  reg        [21:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_5;
  reg        [25:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_4;
  reg        [6:0]    EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_9;
  reg        [26:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_2;
  reg        [10:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_8;
  reg        [26:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_1;
  reg        [26:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_3;
  reg        [30:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0;
  wire       [6:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_9;
  wire       [10:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8;
  wire       [2:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_7;
  wire       [14:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6;
  wire       [21:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5;
  wire       [25:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4;
  wire       [26:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3;
  wire       [26:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2;
  wire       [26:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1;
  wire       [30:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0;
  reg        [3:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_62;
  reg        [6:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_59;
  reg        [7:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_58;
  reg        [1:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_64;
  reg        [2:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_63;
  reg        [0:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_65;
  reg        [4:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_61;
  reg        [13:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_47;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_60;
  reg        [12:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_46;
  reg        [18:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_45;
  reg        [18:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_44;
  reg        [18:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_43;
  reg        [18:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_42;
  reg        [8:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_57;
  reg        [13:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_35;
  reg        [9:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_56;
  reg        [12:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_34;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_33;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_32;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_31;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_30;
  reg        [10:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_55;
  reg        [11:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_29;
  reg        [13:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_25;
  reg        [12:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_24;
  reg        [12:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_53;
  reg        [11:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_23;
  reg        [13:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_52;
  reg        [13:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_21;
  reg        [17:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_48;
  reg        [12:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_20;
  reg        [11:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_41;
  reg        [11:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_19;
  reg        [10:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_40;
  reg        [10:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_18;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_17;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_15;
  reg        [18:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_39;
  reg        [13:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_14;
  reg        [21:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_36;
  reg        [12:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_13;
  reg        [11:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_54;
  reg        [10:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_28;
  reg        [11:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_12;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_27;
  reg        [10:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_11;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_10;
  reg        [14:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_51;
  reg        [19:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_38;
  reg        [20:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_37;
  reg        [23:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_26;
  reg        [15:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_50;
  reg        [10:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_22;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_16;
  reg        [16:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_49;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_9;
  reg        [21:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_8;
  reg        [21:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_6;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_5;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_4;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_3;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_2;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_7;
  reg        [22:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0;
  wire       [0:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_65;
  wire       [1:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_64;
  wire       [2:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_63;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_62;
  wire       [4:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_61;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_60;
  wire       [6:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_59;
  wire       [7:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_58;
  wire       [8:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_57;
  wire       [9:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_56;
  wire       [10:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_55;
  wire       [11:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_54;
  wire       [12:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_53;
  wire       [13:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_52;
  wire       [14:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_51;
  wire       [15:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_50;
  wire       [16:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_49;
  wire       [17:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_48;
  wire       [13:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_47;
  wire       [12:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_46;
  wire       [18:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_45;
  wire       [18:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_44;
  wire       [18:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_43;
  wire       [18:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_42;
  wire       [11:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_41;
  wire       [10:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_40;
  wire       [18:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_39;
  wire       [19:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_38;
  wire       [20:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_37;
  wire       [21:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_36;
  wire       [13:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_35;
  wire       [12:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_34;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_33;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_32;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_31;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_30;
  wire       [11:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_29;
  wire       [10:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_28;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_27;
  wire       [23:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_26;
  wire       [13:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_25;
  wire       [12:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_24;
  wire       [11:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_23;
  wire       [10:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_22;
  wire       [13:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_21;
  wire       [12:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_20;
  wire       [11:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_19;
  wire       [10:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_18;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_17;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_16;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_15;
  wire       [13:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_14;
  wire       [12:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_13;
  wire       [11:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_12;
  wire       [10:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_11;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_10;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_9;
  wire       [21:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7;
  wire       [21:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1;
  wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [0:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_63 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [1:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_61 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [2:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_59 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [3:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_57 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [4:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_55 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [5:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_53 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [6:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_51 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [7:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_49 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [8:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_47 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [9:0]    EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_45 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [10:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_43 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [11:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_41 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [12:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_39 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [13:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_37 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [14:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_35 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [15:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_33 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [16:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_31 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [17:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_29 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [18:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_27 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_25 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [20:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_23 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [21:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_21 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [22:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_19 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [23:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_17 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [24:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_15 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [25:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_13 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [26:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_11 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [27:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_9 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [28:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_7 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [29:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_5 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [30:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [32:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [32:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1 /* synthesis syn_keep = 1 */ ;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_SIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
  wire       [1:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
  wire       [0:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [31:0]   FrontendPlugin_allocated_PC_0;
  reg                 CommitPlugin_logic_commit_continue_1;
  wire       [0:0]    FrontendPlugin_allocated_ROB_MSB_0;
  wire       [1:0]    FrontendPlugin_decompressed_GSHARE_COUNTER_0_0;
  wire       [0:0]    FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_0;
  reg        [6:0]    FetchPlugin_stages_1_GSharePlugin_logic_HASH;
  reg                 FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_valid;
  reg        [6:0]    FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_address;
  reg        [1:0]    FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_0;
  wire                FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_valid;
  wire       [6:0]    FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [23:0]   FetchPlugin_stages_0_BRANCH_HISTORY;
  wire       [6:0]    FetchPlugin_stages_0_GSharePlugin_logic_HASH;
  reg                 _zz_26;
  wire                FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALUE;
  wire                FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALID;
  wire       [31:0]   FetchPlugin_stages_1_Prediction_WORD_BRANCH_PC_NEXT;
  wire                FetchPlugin_stages_1_Prediction_WORD_BRANCH_VALID;
  (* keep , syn_keep *) reg        [1:0]    FetchPlugin_stages_1_GSHARE_COUNTER_0 /* synthesis syn_keep = 1 */ ;
  wire                FetchPlugin_stages_1_BtbPlugin_logic_HIT;
  (* keep , syn_keep *) wire       [15:0]   FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_pcTarget /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_isBranch /* synthesis syn_keep = 1 */ ;
  reg                 _zz_27;
  reg                 _zz_28;
  wire       [3:0]    FrontendPlugin_allocated_ROB_ID /* verilator public */ ;
  reg                 _zz_29;
  wire                FrontendPlugin_allocated_BRANCH_EARLY_0_taken;
  wire       [31:0]   FrontendPlugin_allocated_BRANCH_EARLY_0_pc;
  reg        [2:0]    BranchContextPlugin_logic_alloc_allocNext_1;
  wire                FrontendPlugin_allocated_BRANCH_SEL_0;
  wire       [1:0]    FrontendPlugin_allocated_BRANCH_ID_0;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RD_0;
  wire                FrontendPlugin_allocated_WRITE_RD_0;
  wire                FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0;
  wire                FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_0;
  wire       [31:0]   FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_0;
  wire       [31:0]   FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_0;
  wire                FrontendPlugin_aligned_isFlushed;
  reg        [31:0]   AlignerPlugin_setup_s2m_Fetch_FETCH_PC_INC;
  wire                AlignerPlugin_setup_s2m_isFlushed;
  reg                 AlignerPlugin_setup_s2m_ready;
  wire                FrontendPlugin_aligned_ready;
  reg                 AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE;
  reg                 AlignerPlugin_setup_s2m_Fetch_WORD_FAULT;
  reg                 FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0;
  reg                 FrontendPlugin_aligned_Frontend_FETCH_FAULT_0;
  reg        [11:0]   AlignerPlugin_setup_s2m_FETCH_ID;
  reg        [11:0]   FrontendPlugin_aligned_FETCH_ID_0;
  reg        [31:0]   AlignerPlugin_setup_s2m_Fetch_FETCH_PC;
  reg        [1:0]    AlignerPlugin_setup_s2m_GSHARE_COUNTER_0;
  reg        [1:0]    FrontendPlugin_aligned_GSHARE_COUNTER_0_0;
  reg                 AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE;
  reg                 FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_0;
  reg                 AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID;
  reg                 FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_0;
  reg        [23:0]   AlignerPlugin_setup_s2m_BRANCH_HISTORY;
  reg        [23:0]   FrontendPlugin_aligned_BRANCH_HISTORY_0;
  reg        [31:0]   AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT;
  reg        [31:0]   FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  reg                 FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0;
  wire       [31:0]   FrontendPlugin_aligned_PC_0;
  wire                FrontendPlugin_aligned_Frontend_MASK_ALIGNED_0;
  wire       [31:0]   FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_0;
  reg        [1:0]    AlignerPlugin_logic_slices_remains_1;
  reg        [1:0]    AlignerPlugin_logic_slices_carry_1;
  reg        [1:0]    AlignerPlugin_logic_slices_used_1;
  reg        [0:0]    AlignerPlugin_setup_s2m_MASK_FRONT;
  reg        [31:0]   AlignerPlugin_setup_s2m_Fetch_WORD;
  reg                 AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID;
  reg        [0:0]    AlignerPlugin_setup_s2m_MASK_BACK;
  wire       [0:0]    FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT;
  wire                AlignerPlugin_setup_s2m_isFlushingRoot;
  reg        [23:0]   FetchPlugin_stages_2_BRANCH_HISTORY;
  reg                 FetchPlugin_stages_2_MMU_IO;
  reg        [31:0]   FetchPlugin_stages_2_MMU_TRANSLATED;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HIT;
  reg                 FetchPlugin_stages_2_MMU_REDO;
  wire                FetchPlugin_stages_2_ready;
  reg                 _zz_FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552;
  reg                 _zz_FetchPlugin_stages_2_isFlushingRoot;
  reg                 FetchPlugin_stages_2_MMU_ALLOW_EXECUTE;
  reg                 FetchPlugin_stages_2_MMU_PAGE_FAULT;
  reg                 FetchPlugin_stages_2_MMU_ACCESS_FAULT;
  wire                FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_error;
  reg        [23:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_address;
  wire                FetchPlugin_stages_2_Fetch_WORD_FAULT;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_FETCH_PC;
  wire                FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HIT;
  wire                FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION;
  wire                FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_0;
  wire       [5:0]    FetchPlugin_stages_1_MMU_WAYS_OH;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_error;
  reg        [23:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address;
  reg        [31:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_0;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_0;
  wire       [31:0]   FetchPlugin_stages_2_Fetch_WORD;
  reg        [31:0]   FetchPlugin_stages_1_Fetch_FETCH_PC;
  wire       [31:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_0;
  wire       [31:0]   FetchPlugin_stages_0_Fetch_FETCH_PC;
  reg                 FetchPlugin_stages_0_ready;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_error;
  wire       [23:0]   FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_address;
  wire       [31:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_0;
  reg                 _zz_30;
  reg        [31:0]   PcPlugin_logic_jump_target_1;
  wire                FetchPlugin_stages_1_isFlushed;
  wire                FetchPlugin_stages_1_ready;
  reg        [11:0]   FetchPlugin_stages_1_FETCH_ID /* verilator public */ ;
  reg                 FrontendPlugin_allocated_ready;
  reg                 FrontendPlugin_decoded_ready;
  wire       [11:0]   FrontendPlugin_allocated_FETCH_ID_0 /* verilator public */ ;
  wire       [11:0]   FrontendPlugin_decoded_FETCH_ID_0 /* verilator public */ ;
  reg                 MmuPlugin_setup_cacheLoad_cmd_valid;
  wire                MmuPlugin_setup_cacheLoad_cmd_ready;
  wire       [31:0]   MmuPlugin_setup_cacheLoad_cmd_payload_virtual;
  wire       [1:0]    MmuPlugin_setup_cacheLoad_cmd_payload_size;
  wire                MmuPlugin_setup_cacheLoad_cmd_payload_redoOnDataHazard;
  wire                MmuPlugin_setup_cacheLoad_cmd_payload_unlocked;
  wire                MmuPlugin_setup_cacheLoad_cmd_payload_unique;
  wire       [31:0]   MmuPlugin_setup_cacheLoad_translated_physical;
  wire                MmuPlugin_setup_cacheLoad_translated_abord;
  wire       [2:0]    MmuPlugin_setup_cacheLoad_cancels;
  wire                MmuPlugin_setup_cacheLoad_rsp_valid;
  wire       [31:0]   MmuPlugin_setup_cacheLoad_rsp_payload_data;
  wire                MmuPlugin_setup_cacheLoad_rsp_payload_fault;
  wire                MmuPlugin_setup_cacheLoad_rsp_payload_redo;
  wire       [1:0]    MmuPlugin_setup_cacheLoad_rsp_payload_refillSlot;
  wire                MmuPlugin_setup_cacheLoad_rsp_payload_refillSlotAny;
  reg                 MmuPlugin_setup_invalidatePort_cmd_valid;
  reg                 MmuPlugin_setup_invalidatePort_rsp_valid;
  wire       [31:0]   _zz_FetchPlugin_stages_1_MMU_IO;
  wire                FetchPlugin_stages_0_valid;
  reg                 _zz_FetchPlugin_stages_1_valid;
  reg                 FetchPlugin_stages_1_valid;
  reg                 _zz_FetchPlugin_stages_2_valid;
  reg                 FetchPlugin_stages_2_valid;
  reg                 _zz_AlignerPlugin_setup_s2m_valid;
  wire                FetchCachePlugin_mem_cmd_valid;
  wire                FetchCachePlugin_mem_cmd_ready;
  wire       [31:0]   FetchCachePlugin_mem_cmd_payload_address;
  wire                FetchCachePlugin_mem_cmd_payload_io;
  wire                FetchCachePlugin_mem_rsp_valid;
  wire                FetchCachePlugin_mem_rsp_ready;
  wire       [31:0]   FetchCachePlugin_mem_rsp_payload_data;
  wire                FetchCachePlugin_mem_rsp_payload_error;
  reg                 FetchCachePlugin_setup_redoJump_valid;
  wire       [31:0]   FetchCachePlugin_setup_redoJump_payload_pc;
  wire                FetchCachePlugin_setup_historyJump_valid;
  wire       [23:0]   FetchCachePlugin_setup_historyJump_payload_history;
  reg                 FetchCachePlugin_setup_invalidatePort_cmd_valid;
  reg                 FetchCachePlugin_setup_invalidatePort_rsp_valid;
  wire                AlignerPlugin_setup_s2m_valid;
  wire                AlignerPlugin_setup_sequenceJump_valid;
  wire       [31:0]   AlignerPlugin_setup_sequenceJump_payload_pc;
  wire                AlignerPlugin_setup_singleFetch;
  wire                FrontendPlugin_aligned_valid;
  wire                FrontendPlugin_decompressed_valid;
  wire                FrontendPlugin_decoded_valid;
  reg                 _zz_FrontendPlugin_serialized_valid;
  reg                 FrontendPlugin_serialized_valid;
  wire                FrontendPlugin_allocated_valid;
  reg                 _zz_FrontendPlugin_dispatch_valid;
  reg                 FrontendPlugin_dispatch_valid;
  wire                FrontendPlugin_decoded_isFireing /* verilator public */ ;
  wire                FrontendPlugin_allocated_isFireing /* verilator public */ ;
  wire                FrontendPlugin_isBusy;
  wire                FrontendPlugin_isBusyAfterDecode;
  wire                DecoderPlugin_setup_exceptionPort_valid;
  reg        [3:0]    DecoderPlugin_setup_exceptionPort_payload_cause;
  wire       [31:0]   DecoderPlugin_setup_exceptionPort_payload_epc;
  reg        [31:0]   DecoderPlugin_setup_exceptionPort_payload_tval;
  reg                 DecoderPlugin_setup_trapHalt;
  reg                 DecoderPlugin_setup_trapRaise;
  wire                DecoderPlugin_setup_trapReady;
  wire                DecoderPlugin_setup_debugEnter_0;
  wire                BranchContextPlugin_setup_learnValid;
  wire                DecoderPredictionPlugin_setup_decodeJump_valid;
  wire       [31:0]   DecoderPredictionPlugin_setup_decodeJump_payload_pc;
  wire                DecoderPredictionPlugin_setup_historyPush_flush;
  wire       [0:0]    DecoderPredictionPlugin_setup_historyPush_mask;
  wire       [0:0]    DecoderPredictionPlugin_setup_historyPush_taken;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_2_state;
  wire                BtbPlugin_setup_btbJump_valid;
  wire       [31:0]   BtbPlugin_setup_btbJump_payload_pc;
  wire                BtbPlugin_setup_historyPush_flush;
  wire       [0:0]    BtbPlugin_setup_historyPush_mask;
  wire       [0:0]    BtbPlugin_setup_historyPush_taken;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_0_state;
  reg                 Lsu2Plugin_setup_postCommitBusy;
  reg        [1:0]    Lsu2Plugin_setup_fpuWriteSize;
  reg                 Lsu2Plugin_setup_regfilePorts_0_write_valid;
  reg        [5:0]    Lsu2Plugin_setup_regfilePorts_0_write_address;
  reg        [31:0]   Lsu2Plugin_setup_regfilePorts_0_write_data;
  reg        [3:0]    Lsu2Plugin_setup_regfilePorts_0_write_robId;
  reg                 Lsu2Plugin_setup_cacheLoad_cmd_valid;
  wire                Lsu2Plugin_setup_cacheLoad_cmd_ready;
  reg        [31:0]   Lsu2Plugin_setup_cacheLoad_cmd_payload_virtual;
  reg        [1:0]    Lsu2Plugin_setup_cacheLoad_cmd_payload_size;
  reg                 Lsu2Plugin_setup_cacheLoad_cmd_payload_redoOnDataHazard;
  wire                Lsu2Plugin_setup_cacheLoad_cmd_payload_unlocked;
  reg                 Lsu2Plugin_setup_cacheLoad_cmd_payload_unique;
  reg        [31:0]   Lsu2Plugin_setup_cacheLoad_translated_physical;
  reg                 Lsu2Plugin_setup_cacheLoad_translated_abord;
  wire       [2:0]    Lsu2Plugin_setup_cacheLoad_cancels;
  wire                Lsu2Plugin_setup_cacheLoad_rsp_valid;
  wire       [31:0]   Lsu2Plugin_setup_cacheLoad_rsp_payload_data;
  wire                Lsu2Plugin_setup_cacheLoad_rsp_payload_fault;
  wire                Lsu2Plugin_setup_cacheLoad_rsp_payload_redo;
  wire       [1:0]    Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlot;
  wire                Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlotAny;
  reg                 Lsu2Plugin_setup_cacheStore_cmd_valid;
  wire                Lsu2Plugin_setup_cacheStore_cmd_ready;
  reg        [31:0]   Lsu2Plugin_setup_cacheStore_cmd_payload_address;
  reg        [31:0]   Lsu2Plugin_setup_cacheStore_cmd_payload_data;
  wire       [3:0]    Lsu2Plugin_setup_cacheStore_cmd_payload_mask;
  wire                Lsu2Plugin_setup_cacheStore_cmd_payload_generation;
  reg                 Lsu2Plugin_setup_cacheStore_cmd_payload_io;
  reg                 Lsu2Plugin_setup_cacheStore_cmd_payload_flush;
  wire                Lsu2Plugin_setup_cacheStore_cmd_payload_flushFree;
  reg                 Lsu2Plugin_setup_cacheStore_cmd_payload_prefetch;
  wire                Lsu2Plugin_setup_cacheStore_rsp_valid;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_fault;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_redo;
  wire       [1:0]    Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlot;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlotAny;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_generationKo;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_flush;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_prefetch;
  wire       [31:0]   Lsu2Plugin_setup_cacheStore_rsp_payload_address;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_io;
  reg                 Lsu2Plugin_setup_sharedCompletion_valid;
  wire       [3:0]    Lsu2Plugin_setup_sharedCompletion_payload_id;
  reg                 Lsu2Plugin_setup_sharedTrap_valid;
  reg        [3:0]    Lsu2Plugin_setup_sharedTrap_payload_robId;
  reg                 Lsu2Plugin_setup_sharedTrap_payload_trap;
  wire       [31:0]   Lsu2Plugin_setup_sharedTrap_payload_pcTarget;
  reg        [3:0]    Lsu2Plugin_setup_sharedTrap_payload_cause;
  wire       [31:0]   Lsu2Plugin_setup_sharedTrap_payload_tval;
  wire                Lsu2Plugin_setup_sharedTrap_payload_skipCommit;
  reg        [7:0]    Lsu2Plugin_setup_sharedTrap_payload_reason;
  reg                 Lsu2Plugin_setup_specialTrap_valid;
  wire       [3:0]    Lsu2Plugin_setup_specialTrap_payload_robId;
  wire       [3:0]    Lsu2Plugin_setup_specialTrap_payload_cause;
  wire       [31:0]   Lsu2Plugin_setup_specialTrap_payload_tval;
  wire                Lsu2Plugin_setup_specialTrap_payload_skipCommit;
  wire       [7:0]    Lsu2Plugin_setup_specialTrap_payload_reason;
  reg                 Lsu2Plugin_setup_specialCompletion_valid;
  wire       [3:0]    Lsu2Plugin_setup_specialCompletion_payload_id;
  reg                 Lsu2Plugin_setup_flushPort_cmd_valid;
  reg                 Lsu2Plugin_setup_flushPort_cmd_payload_withFree;
  reg                 Lsu2Plugin_setup_flushPort_rsp_valid;
  wire                DataCachePlugin_setup_writebackBusy;
  wire       [1:0]    DataCachePlugin_setup_refillCompletions;
  reg                 DataCachePlugin_setup_lockPort_valid;
  reg        [31:0]   DataCachePlugin_setup_lockPort_address;
  wire                CommitPlugin_setup_jump_valid;
  wire       [31:0]   CommitPlugin_setup_jump_payload_pc;
  wire       [3:0]    CommitPlugin_setup_robLineMask_line;
  reg        [0:0]    CommitPlugin_setup_robLineMask_mask;
  wire                CommitPlugin_setup_isRobEmpty;
  wire                PrivilegedPlugin_io_int_machine_timer /* verilator public */ ;
  wire                PrivilegedPlugin_io_int_machine_software /* verilator public */ ;
  wire                PrivilegedPlugin_io_int_machine_external /* verilator public */ ;
  wire                PrivilegedPlugin_io_int_supervisor_external /* verilator public */ ;
  wire       [63:0]   PrivilegedPlugin_io_rdtime;
  reg                 PrivilegedPlugin_setup_jump_valid;
  reg        [31:0]   PrivilegedPlugin_setup_jump_payload_pc;
  reg        [1:0]    PrivilegedPlugin_setup_privilege;
  wire                PrivilegedPlugin_setup_withMachinePrivilege;
  wire                PrivilegedPlugin_setup_withSupervisorPrivilege;
  reg                 PrivilegedPlugin_setup_xretAwayFromMachine;
  reg                 PrivilegedPlugin_setup_trapEvent;
  reg                 PrivilegedPlugin_setup_redoTriggered;
  wire                PrivilegedPlugin_setup_setFpDirty;
  wire                PrivilegedPlugin_setup_isFpuEnabled;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_valid;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_valid;
  wire                ALU0_IntAluPlugin_setup_intFormatPort_valid;
  wire       [31:0]   ALU0_IntAluPlugin_setup_intFormatPort_payload;
  wire                ALU0_ShiftPlugin_setup_intFormatPort_valid;
  wire       [31:0]   ALU0_ShiftPlugin_setup_intFormatPort_payload;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_valid;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_valid;
  wire                EU0_MulPlugin_setup_intFormatPort_valid;
  wire       [31:0]   EU0_MulPlugin_setup_intFormatPort_payload;
  wire                EU0_DivPlugin_setup_intFormatPort_valid;
  wire       [31:0]   EU0_DivPlugin_setup_intFormatPort_payload;
  wire                EU0_BranchPlugin_setup_intFormatPort_valid;
  wire       [31:0]   EU0_BranchPlugin_setup_intFormatPort_payload;
  wire                EU0_BranchPlugin_setup_reschedule_valid;
  wire       [3:0]    EU0_BranchPlugin_setup_reschedule_payload_robId;
  wire                EU0_BranchPlugin_setup_reschedule_payload_trap;
  wire       [31:0]   EU0_BranchPlugin_setup_reschedule_payload_pcTarget;
  wire       [3:0]    EU0_BranchPlugin_setup_reschedule_payload_cause;
  wire       [31:0]   EU0_BranchPlugin_setup_reschedule_payload_tval;
  wire                EU0_BranchPlugin_setup_reschedule_payload_skipCommit;
  wire       [7:0]    EU0_BranchPlugin_setup_reschedule_payload_reason;
  wire                AguPlugin_setup_port_valid /* verilator public */ ;
  wire       [3:0]    AguPlugin_setup_port_payload_robId /* verilator public */ ;
  wire       [0:0]    AguPlugin_setup_port_payload_robIdMsb;
  wire       [3:0]    AguPlugin_setup_port_payload_aguId /* verilator public */ ;
  wire                AguPlugin_setup_port_payload_load /* verilator public */ ;
  wire       [31:0]   AguPlugin_setup_port_payload_address;
  wire       [1:0]    AguPlugin_setup_port_payload_size;
  wire                AguPlugin_setup_port_payload_unsigned;
  wire       [5:0]    AguPlugin_setup_port_payload_physicalRd;
  wire                AguPlugin_setup_port_payload_writeRd;
  wire       [31:0]   AguPlugin_setup_port_payload_pc;
  wire                AguPlugin_setup_port_payload_lr;
  wire                AguPlugin_setup_port_payload_earlySample;
  wire       [31:0]   AguPlugin_setup_port_payload_earlyPc;
  wire       [31:0]   AguPlugin_setup_port_payload_data /* verilator public */ ;
  wire                AguPlugin_setup_port_payload_amo;
  wire                AguPlugin_setup_port_payload_sc;
  wire                AguPlugin_setup_port_payload_swap;
  wire       [2:0]    AguPlugin_setup_port_payload_op;
  wire                EnvCallPlugin_setup_reschedule_valid;
  wire       [3:0]    EnvCallPlugin_setup_reschedule_payload_robId;
  reg        [3:0]    EnvCallPlugin_setup_reschedule_payload_cause;
  reg        [31:0]   EnvCallPlugin_setup_reschedule_payload_tval;
  reg                 EnvCallPlugin_setup_reschedule_payload_skipCommit;
  reg        [7:0]    EnvCallPlugin_setup_reschedule_payload_reason;
  wire                EU0_CsrAccessPlugin_setup_intFormatPort_valid;
  wire       [31:0]   EU0_CsrAccessPlugin_setup_intFormatPort_payload;
  reg                 EU0_CsrAccessPlugin_setup_onDecodeTrap;
  reg                 EU0_CsrAccessPlugin_setup_onDecodeFlushPipeline;
  wire                EU0_CsrAccessPlugin_setup_onDecodeRead;
  wire                EU0_CsrAccessPlugin_setup_onDecodeWrite;
  wire       [11:0]   EU0_CsrAccessPlugin_setup_onDecodeAddress;
  reg                 EU0_CsrAccessPlugin_setup_onReadHalt;
  reg                 EU0_CsrAccessPlugin_setup_onWriteHalt;
  reg        [31:0]   EU0_CsrAccessPlugin_setup_onReadToWriteBits;
  reg        [31:0]   EU0_CsrAccessPlugin_setup_onWriteBits;
  wire       [11:0]   EU0_CsrAccessPlugin_setup_onWriteAddress;
  wire                EU0_CsrAccessPlugin_setup_onWriteFlushPipeline;
  wire       [11:0]   EU0_CsrAccessPlugin_setup_onReadAddress;
  wire                EU0_CsrAccessPlugin_setup_onReadMovingOff;
  wire                EU0_CsrAccessPlugin_setup_onWriteMovingOff;
  wire                EU0_CsrAccessPlugin_setup_trap_valid;
  wire       [3:0]    EU0_CsrAccessPlugin_setup_trap_payload_robId;
  reg        [3:0]    EU0_CsrAccessPlugin_setup_trap_payload_cause;
  wire       [31:0]   EU0_CsrAccessPlugin_setup_trap_payload_tval;
  wire                EU0_CsrAccessPlugin_setup_trap_payload_skipCommit;
  wire       [7:0]    EU0_CsrAccessPlugin_setup_trap_payload_reason;
  wire                FetchPlugin_stages_1_isFireing;
  reg                 _zz_FetchPlugin_stages_1_isFirstCycle;
  wire                when_Stage_l170;
  wire                FetchPlugin_stages_1_isFirstCycle /* verilator public */ ;
  wire       [5:0]    _zz_PcPlugin_logic_jump_oh;
  wire                _zz_PcPlugin_logic_jump_oh_1;
  wire                _zz_PcPlugin_logic_jump_oh_2;
  wire                _zz_PcPlugin_logic_jump_oh_3;
  wire                _zz_PcPlugin_logic_jump_oh_4;
  wire                _zz_PcPlugin_logic_jump_oh_5;
  reg        [5:0]    _zz_PcPlugin_logic_jump_oh_6;
  wire                _zz_PcPlugin_logic_jump_oh_7;
  wire       [5:0]    PcPlugin_logic_jump_oh;
  (* keep , syn_keep *) wire       [31:0]   PcPlugin_logic_jump_target /* synthesis syn_keep = 1 */ ;
  wire                _zz_PcPlugin_logic_jump_target_1;
  wire                when_PcPlugin_l57;
  wire                PcPlugin_logic_jump_pcLoad_valid;
  wire       [31:0]   PcPlugin_logic_jump_pcLoad_payload_pc;
  wire                FetchCachePlugin_logic_translationPort_wake;
  wire                FetchCachePlugin_logic_banks_0_write_valid;
  wire       [5:0]    FetchCachePlugin_logic_banks_0_write_payload_address;
  wire       [31:0]   FetchCachePlugin_logic_banks_0_write_payload_data;
  wire                FetchCachePlugin_logic_banks_0_read_cmd_valid;
  wire       [5:0]    FetchCachePlugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [31:0]   FetchCachePlugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [0:0]    FetchCachePlugin_logic_waysWrite_mask;
  reg        [1:0]    FetchCachePlugin_logic_waysWrite_address;
  reg                 FetchCachePlugin_logic_waysWrite_tag_loaded;
  reg                 FetchCachePlugin_logic_waysWrite_tag_error;
  reg        [23:0]   FetchCachePlugin_logic_waysWrite_tag_address;
  wire                FetchCachePlugin_logic_ways_0_read_cmd_valid;
  wire       [1:0]    FetchCachePlugin_logic_ways_0_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_0_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_0_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [23:0]   FetchCachePlugin_logic_ways_0_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [25:0]   _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded;
  reg                 FetchCachePlugin_logic_plru_write_valid;
  reg        [1:0]    FetchCachePlugin_logic_plru_write_payload_address;
  reg                 FetchCachePlugin_logic_invalidate_requested;
  reg                 FetchCachePlugin_logic_invalidate_canStart;
  reg        [2:0]    FetchCachePlugin_logic_invalidate_counter;
  wire                FetchCachePlugin_logic_invalidate_done;
  reg                 FetchCachePlugin_logic_invalidate_firstEver;
  wire                when_FetchCachePlugin_l379;
  wire                when_FetchCachePlugin_l383;
  wire                FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l389;
  wire                when_FetchCachePlugin_l391;
  wire                when_FetchCachePlugin_l396;
  reg                 FetchCachePlugin_logic_invalidate_done_regNext;
  wire                when_FetchCachePlugin_l400;
  reg                 FetchCachePlugin_logic_refill_start_valid;
  wire       [31:0]   FetchCachePlugin_logic_refill_start_address;
  wire                FetchCachePlugin_logic_refill_start_isIo;
  reg                 FetchCachePlugin_logic_refill_fire;
  reg                 FetchCachePlugin_logic_refill_valid;
  (* keep , syn_keep *) reg        [31:0]   FetchCachePlugin_logic_refill_address /* synthesis syn_keep = 1 */ ;
  reg                 FetchCachePlugin_logic_refill_isIo;
  reg                 FetchCachePlugin_logic_refill_hadError;
  reg        [31:0]   FetchCachePlugin_logic_refill_pushCounter;
  wire                when_FetchCachePlugin_l422;
  reg                 FetchCachePlugin_logic_refill_cmdSent;
  wire                FetchCachePlugin_mem_cmd_fire;
  wire                when_Utils_l578;
  reg                 FetchCachePlugin_logic_refill_randomWay_willIncrement;
  wire                FetchCachePlugin_logic_refill_randomWay_willClear;
  wire                FetchCachePlugin_logic_refill_randomWay_willOverflowIfInc;
  wire                FetchCachePlugin_logic_refill_randomWay_willOverflow;
  (* keep , syn_keep *) reg        [3:0]    FetchCachePlugin_logic_refill_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                when_FetchCachePlugin_l470;
  wire                FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l476;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_0;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_1;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_2;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_3;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_4;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_5;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_translatedHits;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_bypassHits;
  reg                 FetchCachePlugin_logic_read_ctrl_redoIt;
  wire                FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552;
  wire                FetchPlugin_stages_2_isFireing;
  wire                when_FetchCachePlugin_l562;
  wire                FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l583;
  wire                when_FetchCachePlugin_l593;
  wire                AlignerPlugin_logic_ignoreInput;
  wire                AlignerPlugin_logic_isInputValid;
  wire                when_AlignerPlugin_l98;
  reg        [31:0]   AlignerPlugin_logic_buffer_data;
  reg        [0:0]    AlignerPlugin_logic_buffer_mask;
  reg        [31:0]   AlignerPlugin_logic_buffer_pc;
  reg                 AlignerPlugin_logic_buffer_fault;
  reg                 AlignerPlugin_logic_buffer_fault_page;
  reg                 AlignerPlugin_logic_buffer_branchValid;
  reg        [31:0]   AlignerPlugin_logic_buffer_branchPcNext;
  reg        [23:0]   AlignerPlugin_logic_buffer_wordContexts_0;
  reg                 AlignerPlugin_logic_buffer_wordContexts_1;
  reg                 AlignerPlugin_logic_buffer_wordContexts_3;
  reg        [1:0]    AlignerPlugin_logic_buffer_wordContexts_4_0;
  reg        [11:0]   AlignerPlugin_logic_buffer_firstWordContexts_0;
  wire       [63:0]   _zz_AlignerPlugin_logic_slices_data_0;
  wire       [31:0]   AlignerPlugin_logic_slices_data_0;
  wire       [31:0]   AlignerPlugin_logic_slices_data_1;
  wire       [1:0]    AlignerPlugin_logic_slices_carry;
  wire       [1:0]    AlignerPlugin_logic_slices_remains;
  wire       [1:0]    AlignerPlugin_logic_slices_used;
  wire       [1:0]    AlignerPlugin_logic_decoders_0_usage;
  wire                AlignerPlugin_logic_decoders_0_notEnoughData;
  wire                AlignerPlugin_logic_decoders_0_pastPrediction;
  wire                AlignerPlugin_logic_decoders_0_usable;
  wire       [1:0]    AlignerPlugin_logic_decoders_1_usage;
  wire                AlignerPlugin_logic_decoders_1_notEnoughData;
  wire                AlignerPlugin_logic_decoders_1_pastPrediction;
  wire                AlignerPlugin_logic_decoders_1_usable;
  wire                _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0;
  wire       [1:0]    _zz_AlignerPlugin_logic_extractors_0_maskOh;
  wire                _zz_AlignerPlugin_logic_extractors_0_maskOh_1;
  reg        [1:0]    _zz_AlignerPlugin_logic_extractors_0_maskOh_2;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_maskOh;
  wire                _zz_AlignerPlugin_logic_extractors_0_usage;
  wire                _zz_AlignerPlugin_logic_extractors_0_usage_1;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_usage;
  wire                AlignerPlugin_logic_extractors_0_usable;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_slice0;
  wire                AlignerPlugin_logic_extractors_0_valid;
  wire                AlignerPlugin_logic_extractors_0_bufferPredictionLast;
  wire                AlignerPlugin_logic_extractors_0_inputPredictionLast;
  wire                AlignerPlugin_logic_extractors_0_lastWord;
  wire                _zz_AlignerPlugin_logic_extractors_0_sliceOffset;
  wire       [0:0]    AlignerPlugin_logic_extractors_0_sliceOffset;
  wire                AlignerPlugin_logic_extractors_0_firstWord;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_pcWord;
  wire                when_AlignerPlugin_l230;
  wire                when_AlignerPlugin_l235;
  wire                FrontendPlugin_aligned_isFireing;
  wire                AlignerPlugin_logic_fireOutput;
  wire                AlignerPlugin_logic_fireInput;
  wire       [0:0]    AlignerPlugin_logic_postMask;
  reg                 AlignerPlugin_logic_correctionSent;
  wire                when_AlignerPlugin_l264;
  wire                _zz_FetchPlugin_stages_1_isFlushingRoot;
  wire                AlignerPlugin_setup_s2m_haltRequest_AlignerPlugin_l270;
  wire                integer_RfAllocationPlugin_logic_pop_blocked;
  wire                FrontendPlugin_allocated_haltRequest_RfAllocationPlugin_l55;
  wire                when_RfAllocationPlugin_l63;
  reg        [2:0]    BranchContextPlugin_logic_ptr_alloc;
  reg        [2:0]    BranchContextPlugin_logic_ptr_commited;
  reg        [2:0]    BranchContextPlugin_logic_ptr_free;
  wire       [2:0]    BranchContextPlugin_logic_ptr_occupancy;
  wire       [2:0]    BranchContextPlugin_logic_alloc_allocNext;
  reg                 BranchContextPlugin_logic_alloc_full;
  wire                when_BranchContextPlugin_l97;
  wire                when_BranchContextPlugin_l110;
  wire                FrontendPlugin_allocated_haltRequest_BranchContextPlugin_l111;
  reg        [23:0]   HistoryPlugin_logic_onCommit_value /* verilator public */ ;
  wire       [23:0]   HistoryPlugin_logic_onCommit_whitebox_0 /* verilator public */ ;
  reg        [3:0]    DecoderPredictionPlugin_logic_ras_ptr_push;
  reg        [3:0]    DecoderPredictionPlugin_logic_ras_ptr_pop;
  reg                 DecoderPredictionPlugin_logic_ras_ptr_pushIt;
  reg                 DecoderPredictionPlugin_logic_ras_ptr_popIt;
  wire       [31:0]   DecoderPredictionPlugin_logic_ras_read;
  wire                DecoderPredictionPlugin_logic_ras_write_valid;
  wire       [3:0]    DecoderPredictionPlugin_logic_ras_write_payload_address;
  reg        [31:0]   DecoderPredictionPlugin_logic_ras_write_payload_data;
  wire       [31:0]   BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice;
  wire       [31:0]   BranchContextPlugin_learn_BRANCH_FINAL_pcTarget;
  wire                BranchContextPlugin_learn_BRANCH_FINAL_taken;
  wire       [15:0]   BtbPlugin_logic_onLearn_hash;
  wire                BtbPlugin_logic_onLearn_port_valid;
  wire       [2:0]    BtbPlugin_logic_onLearn_port_payload_address;
  wire       [15:0]   BtbPlugin_logic_onLearn_port_payload_data_hash;
  wire       [31:0]   BtbPlugin_logic_onLearn_port_payload_data_pcTarget;
  wire                BtbPlugin_logic_onLearn_port_payload_data_isBranch;
  wire                BranchContextPlugin_free_learn_Prediction_IS_BRANCH;
  wire       [2:0]    BtbPlugin_logic_readCmd_entryAddress;
  wire       [48:0]   _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash;
  wire                BtbPlugin_logic_hitCalc_postPcPrediction;
  wire                BtbPlugin_logic_applyIt_prediction;
  wire                BtbPlugin_logic_applyIt_needIt;
  reg                 BtbPlugin_logic_applyIt_correctionSent;
  wire                when_BtbPlugin_l109;
  wire                BtbPlugin_logic_applyIt_doIt;
  wire                GSharePlugin_logic_mem_write_valid;
  wire       [6:0]    GSharePlugin_logic_mem_write_payload_address;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_0;
  wire       [6:0]    _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH;
  wire                when_GSharePlugin_l98;
  wire       [23:0]   BranchContextPlugin_free_learn_BRANCH_HISTORY;
  wire       [6:0]    _zz_GSharePlugin_logic_onLearn_hash;
  wire       [6:0]    GSharePlugin_logic_onLearn_hash;
  wire       [1:0]    BranchContextPlugin_free_learn_GSHARE_COUNTER_0;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_0;
  wire       [1:0]    GSharePlugin_logic_onLearn_incrValue;
  reg                 GSharePlugin_logic_onLearn_overflow;
  wire                when_GSharePlugin_l123;
  wire                LsuPlugin_peripheralBus_cmd_valid /* verilator public */ ;
  reg                 LsuPlugin_peripheralBus_cmd_ready /* verilator public */ ;
  wire                LsuPlugin_peripheralBus_cmd_payload_write /* verilator public */ ;
  wire       [31:0]   LsuPlugin_peripheralBus_cmd_payload_address /* verilator public */ ;
  wire       [31:0]   LsuPlugin_peripheralBus_cmd_payload_data /* verilator public */ ;
  wire       [3:0]    LsuPlugin_peripheralBus_cmd_payload_mask /* verilator public */ ;
  wire       [1:0]    LsuPlugin_peripheralBus_cmd_payload_size /* verilator public */ ;
  wire                LsuPlugin_peripheralBus_rsp_valid /* verilator public */ ;
  wire                LsuPlugin_peripheralBus_rsp_payload_error /* verilator public */ ;
  wire       [31:0]   LsuPlugin_peripheralBus_rsp_payload_data /* verilator public */ ;
  wire       [1:0]    DataCachePlugin_logic_load_hits;
  wire                DataCachePlugin_logic_load_hit;
  wire       [1:0]    _zz_DataCachePlugin_logic_load_hits_bools_0;
  wire                DataCachePlugin_logic_load_hits_bools_0;
  wire                DataCachePlugin_logic_load_hits_bools_1;
  reg        [1:0]    _zz_DataCachePlugin_logic_load_oh;
  wire       [1:0]    DataCachePlugin_logic_load_oh;
  wire       [1:0]    DataCachePlugin_logic_load_ohHistory_0;
  wire       [1:0]    DataCachePlugin_logic_load_ohHistory_1;
  wire       [1:0]    DataCachePlugin_logic_load_ohHistory_2;
  wire       [1:0]    _zz_DataCachePlugin_logic_load_ohHistory_0;
  reg        [1:0]    _zz_DataCachePlugin_logic_load_ohHistory_1;
  reg        [1:0]    _zz_DataCachePlugin_logic_load_ohHistory_2;
  wire                _zz_MmuPlugin_setup_cacheLoad_cmd_ready;
  wire                _zz_io_load_translated_physical;
  wire                DataCachePlugin_mem_read_cmd_valid;
  wire                DataCachePlugin_mem_read_cmd_ready;
  wire       [0:0]    DataCachePlugin_mem_read_cmd_payload_id;
  wire       [31:0]   DataCachePlugin_mem_read_cmd_payload_address;
  wire                DataCachePlugin_mem_read_rsp_valid;
  wire                DataCachePlugin_mem_read_rsp_ready;
  wire       [0:0]    DataCachePlugin_mem_read_rsp_payload_id;
  wire       [31:0]   DataCachePlugin_mem_read_rsp_payload_data;
  wire                DataCachePlugin_mem_read_rsp_payload_error;
  wire                DataCachePlugin_mem_write_cmd_valid;
  reg                 DataCachePlugin_mem_write_cmd_ready;
  wire                DataCachePlugin_mem_write_cmd_payload_last;
  wire       [31:0]   DataCachePlugin_mem_write_cmd_payload_fragment_address;
  wire       [31:0]   DataCachePlugin_mem_write_cmd_payload_fragment_data;
  wire       [0:0]    DataCachePlugin_mem_write_cmd_payload_fragment_id;
  wire                DataCachePlugin_mem_write_rsp_valid;
  wire                DataCachePlugin_mem_write_rsp_payload_error;
  wire       [0:0]    DataCachePlugin_mem_write_rsp_payload_id;
  reg        [4:0]    CommitPlugin_logic_ptr_alloc;
  reg        [4:0]    CommitPlugin_logic_ptr_commit;
  reg        [4:0]    CommitPlugin_logic_ptr_free;
  wire       [4:0]    CommitPlugin_logic_ptr_commitRow;
  reg        [4:0]    CommitPlugin_logic_ptr_commitNext;
  wire       [4:0]    CommitPlugin_logic_ptr_allocNext;
  wire                CommitPlugin_logic_ptr_full;
  reg                 CommitPlugin_logic_ptr_empty;
  wire                CommitPlugin_logic_ptr_canFree;
  reg        [0:0]    CommitPlugin_logic_ptr_robLineMaskRsp;
  wire                FrontendPlugin_allocated_haltRequest_CommitPlugin_l95;
  reg                 CommitPlugin_logic_reschedule_fresh;
  reg                 CommitPlugin_logic_reschedule_valid;
  reg                 CommitPlugin_logic_reschedule_trap;
  reg                 CommitPlugin_logic_reschedule_skipCommit;
  reg        [3:0]    CommitPlugin_logic_reschedule_robId;
  reg        [31:0]   CommitPlugin_logic_reschedule_pcTarget;
  reg        [3:0]    CommitPlugin_logic_reschedule_cause;
  reg        [31:0]   CommitPlugin_logic_reschedule_tval;
  reg        [7:0]    CommitPlugin_logic_reschedule_reason;
  wire       [3:0]    CommitPlugin_logic_reschedule_commit_row;
  wire                CommitPlugin_logic_reschedule_commit_rowHit;
  wire       [3:0]    CommitPlugin_logic_reschedule_age;
  wire       [3:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_0_age;
  wire       [3:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_1_age;
  wire       [3:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_2_age;
  wire       [3:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_3_age;
  wire       [3:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_4_age;
  reg        [4:0]    CommitPlugin_logic_reschedule_portsLogic_hits;
  wire                when_CommitPlugin_l131;
  wire                _zz_CommitPlugin_logic_reschedule_trap;
  wire                _zz_CommitPlugin_logic_reschedule_trap_1;
  wire                _zz_CommitPlugin_logic_reschedule_trap_2;
  wire                _zz_CommitPlugin_logic_reschedule_trap_3;
  wire                _zz_CommitPlugin_logic_reschedule_trap_4;
  wire                CommitPlugin_logic_reschedule_reschedulePort_valid;
  wire       [3:0]    CommitPlugin_logic_reschedule_reschedulePort_payload_robId;
  wire                CommitPlugin_logic_reschedule_reschedulePort_payload_trap;
  wire       [3:0]    CommitPlugin_logic_reschedule_reschedulePort_payload_cause;
  wire       [31:0]   CommitPlugin_logic_reschedule_reschedulePort_payload_tval;
  wire       [7:0]    CommitPlugin_logic_reschedule_reschedulePort_payload_reason;
  wire                CommitPlugin_logic_reschedule_reschedulePort_payload_skipCommit;
  reg                 CommitPlugin_logic_commit_rescheduleHit;
  wire       [0:0]    CommitPlugin_logic_commit_active;
  reg        [0:0]    CommitPlugin_logic_commit_mask;
  reg        [0:0]    CommitPlugin_logic_commit_maskComb;
  wire                CommitPlugin_logic_commit_lineCommited;
  wire       [3:0]    CommitPlugin_logic_commit_event_robId;
  reg        [0:0]    CommitPlugin_logic_commit_event_mask;
  reg                 CommitPlugin_logic_commit_lineEvent_valid;
  wire       [3:0]    CommitPlugin_logic_commit_lineEvent_payload_robId;
  wire       [0:0]    CommitPlugin_logic_commit_lineEvent_payload_mask;
  wire                CommitPlugin_logic_commit_reschedulePort_valid;
  wire       [3:0]    CommitPlugin_logic_commit_reschedulePort_payload_robId;
  wire       [3:0]    CommitPlugin_logic_commit_reschedulePort_payload_robIdNext;
  wire                CommitPlugin_logic_commit_reschedulePort_payload_trap;
  wire       [3:0]    CommitPlugin_logic_commit_reschedulePort_payload_cause;
  wire       [31:0]   CommitPlugin_logic_commit_reschedulePort_payload_tval;
  wire       [7:0]    CommitPlugin_logic_commit_reschedulePort_payload_reason;
  wire                CommitPlugin_logic_commit_reschedulePort_payload_skipCommit;
  wire       [3:0]    CommitPlugin_logic_commit_head;
  reg        [3:0]    CommitPlugin_logic_commit_headNext;
  wire                CommitPlugin_logic_commit_continue;
  wire                when_CommitPlugin_l194;
  wire                CommitPlugin_commit_slot_0_enable;
  wire                CommitPlugin_commit_slot_0_readyForCommit;
  wire                CommitPlugin_commit_slot_0_rescheduleHitSlot;
  wire                when_CommitPlugin_l203;
  wire                when_CommitPlugin_l207;
  wire                when_CommitPlugin_l211;
  wire                when_CommitPlugin_l217;
  wire                CommitPlugin_logic_free_lineEventStream_valid;
  wire                CommitPlugin_logic_free_lineEventStream_ready;
  wire       [3:0]    CommitPlugin_logic_free_lineEventStream_payload_robId;
  wire       [0:0]    CommitPlugin_logic_free_lineEventStream_payload_mask;
  wire                CommitPlugin_logic_free_robHit;
  wire                CommitPlugin_logic_free_hit;
  wire                CommitPlugin_logic_free_port_valid;
  wire       [3:0]    CommitPlugin_logic_free_port_payload_robId;
  wire       [0:0]    CommitPlugin_logic_free_port_payload_commited;
  wire                robToPc_valid /* verilator public */ ;
  wire       [3:0]    robToPc_robId /* verilator public */ ;
  wire       [31:0]   robToPc_pc_0 /* verilator public */ ;
  wire       [3:0]    commit_robId /* verilator public */ ;
  wire       [0:0]    commit_mask /* verilator public */ ;
  wire                reschedule_valid /* verilator public */ ;
  wire       [3:0]    reschedule_payload_robId /* verilator public */ ;
  wire       [3:0]    reschedule_payload_robIdNext /* verilator public */ ;
  wire                reschedule_payload_trap /* verilator public */ ;
  wire       [3:0]    reschedule_payload_cause /* verilator public */ ;
  wire       [31:0]   reschedule_payload_tval /* verilator public */ ;
  wire       [7:0]    reschedule_payload_reason /* verilator public */ ;
  wire                reschedule_payload_skipCommit /* verilator public */ ;
  wire       [7:0]    rescheduleReason /* verilator public */ ;
  wire       [31:0]   commit_pc_0 /* verilator public */ ;
  wire       [16:0]   CommitDebugFilterPlugin_logic_commits;
  reg        [31:0]   CommitDebugFilterPlugin_logic_filters_0_value;
  reg        [31:0]   CommitDebugFilterPlugin_logic_filters_1_value;
  reg        [31:0]   CommitDebugFilterPlugin_logic_filters_2_value;
  wire       [1:0]    PrivilegedPlugin_logic_defaultTrap_csrPrivilege;
  wire                PrivilegedPlugin_logic_defaultTrap_csrReadOnly;
  wire                when_PrivilegedPlugin_l165;
  reg                 PrivilegedPlugin_logic_machine_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_machine_cause_code;
  reg                 PrivilegedPlugin_logic_machine_mstatus_mie;
  reg                 PrivilegedPlugin_logic_machine_mstatus_mpie;
  reg        [1:0]    PrivilegedPlugin_logic_machine_mstatus_mpp;
  reg        [1:0]    PrivilegedPlugin_logic_machine_mstatus_fs;
  reg                 PrivilegedPlugin_logic_machine_mstatus_sd;
  wire                when_PrivilegedPlugin_l393;
  reg                 PrivilegedPlugin_logic_machine_mstatus_tsr;
  reg                 PrivilegedPlugin_logic_machine_mstatus_tvm;
  reg                 PrivilegedPlugin_logic_machine_mstatus_tw;
  reg                 PrivilegedPlugin_logic_machine_mip_meip;
  reg                 PrivilegedPlugin_logic_machine_mip_mtip;
  reg                 PrivilegedPlugin_logic_machine_mip_msip;
  reg                 PrivilegedPlugin_logic_machine_mie_meie;
  reg                 PrivilegedPlugin_logic_machine_mie_mtie;
  reg                 PrivilegedPlugin_logic_machine_mie_msie;
  reg                 PrivilegedPlugin_logic_machine_medeleg_iam;
  reg                 PrivilegedPlugin_logic_machine_medeleg_bp;
  reg                 PrivilegedPlugin_logic_machine_medeleg_eu;
  reg                 PrivilegedPlugin_logic_machine_medeleg_es;
  reg                 PrivilegedPlugin_logic_machine_medeleg_ipf;
  reg                 PrivilegedPlugin_logic_machine_medeleg_lpf;
  reg                 PrivilegedPlugin_logic_machine_medeleg_spf;
  reg                 PrivilegedPlugin_logic_machine_mideleg_st;
  reg                 PrivilegedPlugin_logic_machine_mideleg_se;
  reg                 PrivilegedPlugin_logic_machine_mideleg_ss;
  reg                 PrivilegedPlugin_logic_supervisor_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_supervisor_cause_code;
  reg                 PrivilegedPlugin_logic_supervisor_sstatus_sie;
  reg                 PrivilegedPlugin_logic_supervisor_sstatus_spie;
  reg        [0:0]    PrivilegedPlugin_logic_supervisor_sstatus_spp;
  reg                 PrivilegedPlugin_logic_supervisor_sip_seipSoft;
  reg                 PrivilegedPlugin_logic_supervisor_sip_seipInput;
  wire                PrivilegedPlugin_logic_supervisor_sip_seipOr;
  reg                 PrivilegedPlugin_logic_supervisor_sip_stip;
  reg                 PrivilegedPlugin_logic_supervisor_sip_ssip;
  wire                PrivilegedPlugin_logic_supervisor_sip_seipMasked;
  wire                PrivilegedPlugin_logic_supervisor_sip_stipMasked;
  wire                PrivilegedPlugin_logic_supervisor_sip_ssipMasked;
  reg                 PrivilegedPlugin_logic_supervisor_sie_seie;
  reg                 PrivilegedPlugin_logic_supervisor_sie_stie;
  reg                 PrivilegedPlugin_logic_supervisor_sie_ssie;
  wire                _zz_when_PrivilegedPlugin_l644;
  wire                _zz_when_PrivilegedPlugin_l644_1;
  wire                _zz_when_PrivilegedPlugin_l644_2;
  reg                 PrivilegedPlugin_logic_rescheduleUnbuffered_valid;
  reg                 PrivilegedPlugin_logic_rescheduleUnbuffered_ready;
  reg        [3:0]    PrivilegedPlugin_logic_rescheduleUnbuffered_payload_cause;
  reg        [31:0]   PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc;
  reg        [31:0]   PrivilegedPlugin_logic_rescheduleUnbuffered_payload_tval;
  wire                PrivilegedPlugin_logic_rescheduleUnbuffered_payload_fromCommit;
  wire                PrivilegedPlugin_logic_reschedule_valid;
  reg                 PrivilegedPlugin_logic_reschedule_ready;
  wire       [3:0]    PrivilegedPlugin_logic_reschedule_payload_cause;
  wire       [31:0]   PrivilegedPlugin_logic_reschedule_payload_epc;
  wire       [31:0]   PrivilegedPlugin_logic_reschedule_payload_tval;
  wire                PrivilegedPlugin_logic_reschedule_payload_fromCommit;
  reg                 PrivilegedPlugin_logic_rescheduleUnbuffered_rValid;
  reg        [3:0]    PrivilegedPlugin_logic_rescheduleUnbuffered_rData_cause;
  reg        [31:0]   PrivilegedPlugin_logic_rescheduleUnbuffered_rData_epc;
  reg        [31:0]   PrivilegedPlugin_logic_rescheduleUnbuffered_rData_tval;
  reg                 PrivilegedPlugin_logic_rescheduleUnbuffered_rData_fromCommit;
  wire                when_Stream_l369;
  wire                when_PrivilegedPlugin_l592;
  wire                PrivilegedPlugin_logic_targetMachine;
  reg        [31:0]   PrivilegedPlugin_logic_readed;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_valid;
  wire                ALU0_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   ALU0_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [1:0]    ALU0_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   ALU0_IntFormatPlugin_logic_stages_0_raw;
  reg        [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  reg        [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  reg        [31:0]   ALU0_SrcPlugin_logic_addsub_rs2Patched;
  reg        [31:0]   ALU0_IntAluPlugin_logic_process_bitwise;
  reg        [31:0]   ALU0_IntAluPlugin_logic_process_result;
  wire       [4:0]    ALU0_ShiftPlugin_logic_process_amplitude;
  wire       [31:0]   ALU0_ShiftPlugin_logic_process_reversed;
  wire       [31:0]   ALU0_ShiftPlugin_logic_process_shifted;
  wire       [31:0]   ALU0_ShiftPlugin_logic_process_patched;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_valid;
  wire                EU0_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   EU0_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [3:0]    EU0_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   EU0_IntFormatPlugin_logic_stages_0_raw;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_valid;
  reg                 _zz_EU0_ExecutionUnitBase_pipeline_execute_1_valid;
  reg        [31:0]   EU0_SrcPlugin_logic_addsub_rs2Patched;
  wire                EU0_MulPlugin_logic_wake_wakeRobsSel;
  wire                EU0_MulPlugin_logic_wake_wakeRegFileSel;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_1;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_2;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_3;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_1;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_2;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_3;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_1;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_2;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_3;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_1;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_2;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_3;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_1;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_2;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_3;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_1;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_2;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_3;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_1;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_2;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_3;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_1;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_2;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_3;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_1;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_2;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_3;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_9;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_10;
  reg        [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_11;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_12;
  reg        [12:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_13;
  reg        [13:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_14;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_15;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_16;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_17;
  reg        [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_18;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_19;
  reg        [12:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_20;
  reg        [13:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_21;
  reg        [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_22;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_23;
  reg        [12:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_24;
  reg        [13:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_25;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_26;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_27;
  reg        [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_28;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_29;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_30;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_31;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_32;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_33;
  reg        [12:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_34;
  reg        [13:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_35;
  reg        [21:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_36;
  reg        [20:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_37;
  reg        [19:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_38;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_39;
  reg        [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_40;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_41;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_42;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_43;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_44;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_45;
  reg        [12:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_46;
  reg        [13:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_47;
  reg        [17:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_48;
  reg        [16:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_49;
  reg        [15:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_50;
  reg        [14:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_51;
  reg        [13:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_52;
  reg        [12:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_53;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_54;
  reg        [10:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_55;
  reg        [9:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_56;
  reg        [8:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_57;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_58;
  reg        [6:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_59;
  reg        [5:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_60;
  reg        [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_61;
  reg        [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_62;
  reg        [2:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_63;
  reg        [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_64;
  reg        [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_65;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_valid;
  reg                 _zz_EU0_ExecutionUnitBase_pipeline_execute_2_valid;
  reg        [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0;
  reg        [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_1;
  reg        [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_2;
  reg        [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_3;
  reg        [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_4;
  reg        [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_5;
  reg        [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_6;
  reg        [27:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_7;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_1;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_2;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_3;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_4;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_5;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_6;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_7;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_1;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_2;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_3;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_4;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_5;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_6;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_7;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_1;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_2;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_3;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_4;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_5;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_6;
  reg        [23:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_7;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_1;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_2;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_3;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_4;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_5;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_6;
  reg        [22:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_7;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_1;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_2;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_3;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_4;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_5;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_6;
  reg        [18:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_7;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_1;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_2;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_3;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_4;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_5;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_6;
  reg        [11:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_7;
  reg        [2:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_7;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_1;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_2;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_3;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_4;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_5;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_6;
  reg        [7:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_7;
  reg        [6:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_9;
  reg        [66:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0;
  reg        [66:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_1;
  reg        [66:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_2;
  reg        [66:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_3;
  reg        [66:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_4;
  reg        [66:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_5;
  reg        [66:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_6;
  wire                EU0_DivPlugin_logic_wake_wakeRobsSel;
  wire                EU0_DivPlugin_logic_wake_wakeRegFileSel;
  reg                 EU0_DivPlugin_logic_feed_cmdSent;
  wire                toplevel_EU0_DivPlugin_logic_div_io_cmd_fire;
  wire                when_DivPlugin_l76;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_haltRequest_DivPlugin_l83;
  wire                EU0_ExecutionUnitBase_pipeline_execute_1_haltRequest_DivPlugin_l91;
  wire       [34:0]   EU0_DivPlugin_logic_rsp_selected;
  wire       [34:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT;
  wire                EU0_BranchPlugin_logic_wake_wakeRobsSel;
  wire                EU0_BranchPlugin_logic_wake_wakeRegFileSel;
  wire       [2:0]    switch_Misc_l241;
  reg                 _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
  reg                 _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1;
  reg        [31:0]   EU0_BranchPlugin_logic_process_target_a;
  reg        [31:0]   EU0_BranchPlugin_logic_process_target_b;
  wire       [1:0]    EU0_BranchPlugin_logic_process_slices;
  wire       [2:0]    AguPlugin_logic_func3;
  reg                 AguPlugin_logic_fired;
  wire                when_AguPlugin_l89;
  wire                EU0_CsrAccessPlugin_logic_wake_wakeRobsSel;
  wire                EU0_CsrAccessPlugin_logic_wake_wakeRegFileSel;
  wire                LsuPlugin_peripheralBus_toAxiLite4_a_valid;
  wire                LsuPlugin_peripheralBus_toAxiLite4_a_ready;
  wire                LsuPlugin_peripheralBus_toAxiLite4_a_payload_write;
  wire       [31:0]   LsuPlugin_peripheralBus_toAxiLite4_a_payload_address;
  wire       [31:0]   LsuPlugin_peripheralBus_toAxiLite4_a_payload_data;
  wire       [3:0]    LsuPlugin_peripheralBus_toAxiLite4_a_payload_mask;
  wire       [1:0]    LsuPlugin_peripheralBus_toAxiLite4_a_payload_size;
  wire                LsuPlugin_peripheralBus_toAxiLite4_wRaw_valid;
  reg                 LsuPlugin_peripheralBus_toAxiLite4_wRaw_ready;
  wire                LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_write;
  wire       [31:0]   LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_address;
  wire       [31:0]   LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_data;
  wire       [3:0]    LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_mask;
  wire       [1:0]    LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_size;
  reg                 LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_0;
  reg                 LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_1;
  wire                when_Stream_l1058;
  wire                when_Stream_l1058_1;
  wire                LsuPlugin_peripheralBus_toAxiLite4_a_fire;
  wire                LsuPlugin_peripheralBus_toAxiLite4_wRaw_fire;
  wire                when_Stream_l439;
  reg                 LsuPlugin_peripheralBus_toAxiLite4_w_valid;
  wire                LsuPlugin_peripheralBus_toAxiLite4_w_ready;
  wire                LsuPlugin_peripheralBus_toAxiLite4_w_payload_write;
  wire       [31:0]   LsuPlugin_peripheralBus_toAxiLite4_w_payload_address;
  wire       [31:0]   LsuPlugin_peripheralBus_toAxiLite4_w_payload_data;
  wire       [3:0]    LsuPlugin_peripheralBus_toAxiLite4_w_payload_mask;
  wire       [1:0]    LsuPlugin_peripheralBus_toAxiLite4_w_payload_size;
  reg                 LsuPlugin_peripheralBus_toAxiLite4_writeSel;
  wire       [31:0]   LsuPlugin_peripheralBus_toAxiLite4_addr;
  wire                DataCachePlugin_mem_toAxi4_awRaw_valid;
  reg                 DataCachePlugin_mem_toAxi4_awRaw_ready;
  wire                DataCachePlugin_mem_toAxi4_awRaw_payload_last;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_address;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_data;
  wire       [0:0]    DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_id;
  wire                DataCachePlugin_mem_toAxi4_wRaw_valid;
  wire                DataCachePlugin_mem_toAxi4_wRaw_ready;
  wire                DataCachePlugin_mem_toAxi4_wRaw_payload_last;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_address;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_data;
  wire       [0:0]    DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_id;
  reg                 DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_0;
  reg                 DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_1;
  wire                when_Stream_l1058_2;
  wire                when_Stream_l1058_3;
  wire                DataCachePlugin_mem_toAxi4_awRaw_fire;
  wire                DataCachePlugin_mem_toAxi4_wRaw_fire;
  reg                 DataCachePlugin_mem_toAxi4_awRaw_payload_first;
  wire                when_Stream_l439_1;
  reg                 DataCachePlugin_mem_toAxi4_awFiltred_valid;
  reg                 DataCachePlugin_mem_toAxi4_awFiltred_ready;
  wire                DataCachePlugin_mem_toAxi4_awFiltred_payload_last;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_address;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_data;
  wire       [0:0]    DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_id;
  wire                DataCachePlugin_mem_toAxi4_aw_valid;
  wire                DataCachePlugin_mem_toAxi4_aw_ready;
  wire                DataCachePlugin_mem_toAxi4_aw_payload_last;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_aw_payload_fragment_address;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_aw_payload_fragment_data;
  wire       [0:0]    DataCachePlugin_mem_toAxi4_aw_payload_fragment_id;
  reg                 DataCachePlugin_mem_toAxi4_awFiltred_rValid;
  reg                 DataCachePlugin_mem_toAxi4_awFiltred_rData_last;
  reg        [31:0]   DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_address;
  reg        [31:0]   DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_data;
  reg        [0:0]    DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_id;
  wire                when_Stream_l369_1;
  wire                _zz_DataCachePlugin_mem_toAxi4_wRaw_ready;
  wire                DataCachePlugin_mem_toAxi4_w_valid;
  wire                DataCachePlugin_mem_toAxi4_w_ready;
  wire                DataCachePlugin_mem_toAxi4_w_payload_last;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_w_payload_fragment_address;
  wire       [31:0]   DataCachePlugin_mem_toAxi4_w_payload_fragment_data;
  wire       [0:0]    DataCachePlugin_mem_toAxi4_w_payload_fragment_id;
  wire                FrontendPlugin_allocated_haltRequest_FrontendPlugin_l67;
  wire                integer_RfTranslationPlugin_logic_onCommit_writeRd_0;
  wire       [5:0]    integer_RfTranslationPlugin_logic_onCommit_physRd_0;
  wire       [4:0]    integer_RfTranslationPlugin_logic_onCommit_archRd_0;
  reg        [5:0]    integer_RfTranslationPlugin_logic_init_counter;
  wire                integer_RfTranslationPlugin_logic_init_busy;
  wire                when_RfTranslationPlugin_l193;
  wire                integer_RfAllocationPlugin_logic_push_mask_0;
  wire                integer_RfAllocationPlugin_logic_push_writeRd_0;
  wire       [5:0]    integer_RfAllocationPlugin_logic_push_physicalRdNew_0;
  wire       [5:0]    integer_RfAllocationPlugin_logic_push_physicalRdOld_0;
  wire                when_RfAllocationPlugin_l81;
  reg        [6:0]    integer_RfAllocationPlugin_logic_init_counter;
  wire                integer_RfAllocationPlugin_logic_init_busy;
  wire                BranchContextPlugin_logic_onCommit_isBranch_0;
  wire                BranchContextPlugin_logic_onCommit_isBranchCommit_0;
  wire       [2:0]    BranchContextPlugin_logic_onCommit_commitedNext;
  wire                HistoryPlugin_logic_onCommit_isConditionalBranch_0;
  wire                HistoryPlugin_logic_onCommit_isTaken_0;
  wire       [23:0]   HistoryPlugin_logic_onCommit_valueNext;
  wire                when_HistoryPlugin_l90;
  reg        [23:0]   HistoryPlugin_logic_onFetch_value;
  reg        [23:0]   HistoryPlugin_logic_onFetch_valueNext;
  wire       [23:0]   HistoryPlugin_logic_update_pushes_0_stateNext;
  wire                when_HistoryPlugin_l115;
  wire       [23:0]   HistoryPlugin_logic_update_pushes_2_stateNext;
  wire                when_HistoryPlugin_l115_1;
  wire       [23:0]   HistoryPlugin_logic_update_rescheduleFlush_instHistory;
  wire                HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch;
  wire                HistoryPlugin_logic_update_rescheduleFlush_isTaken;
  wire       [23:0]   HistoryPlugin_logic_update_rescheduleFlush_newHistory;
  wire       [3:0]    DecoderPredictionPlugin_logic_ras_healPush;
  wire       [3:0]    DecoderPredictionPlugin_logic_ras_healPop;
  wire                DecoderPredictionPlugin_logic_decodePatch_rasPushUsed;
  wire                Lsu2Plugin_logic_translationWake;
  wire                Lsu2Plugin_logic_sqWritebackEvent_valid;
  wire       [2:0]    Lsu2Plugin_logic_sqWritebackEvent_payload;
  wire                Lsu2Plugin_logic_sqFeedEvent_valid;
  wire       [2:0]    Lsu2Plugin_logic_sqFeedEvent_payload;
  reg                 Lsu2Plugin_logic_lq_regs_0_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_0_valid;
  reg                 Lsu2Plugin_logic_lq_regs_0_redo;
  reg                 Lsu2Plugin_logic_lq_regs_0_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_0_delete;
  reg                 Lsu2Plugin_logic_lq_regs_0_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_0_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_0_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_0_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed;
  reg        [2:0]    Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315;
  wire                when_Lsu2Plugin_l338;
  reg                 Lsu2Plugin_logic_lq_regs_1_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_1_valid;
  reg                 Lsu2Plugin_logic_lq_regs_1_redo;
  reg                 Lsu2Plugin_logic_lq_regs_1_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_1_delete;
  reg                 Lsu2Plugin_logic_lq_regs_1_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_1_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_1_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_1_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed;
  reg        [2:0]    Lsu2Plugin_logic_lq_regs_1_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_1;
  wire                when_Lsu2Plugin_l338_1;
  reg                 Lsu2Plugin_logic_lq_regs_2_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_2_valid;
  reg                 Lsu2Plugin_logic_lq_regs_2_redo;
  reg                 Lsu2Plugin_logic_lq_regs_2_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_2_delete;
  reg                 Lsu2Plugin_logic_lq_regs_2_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_2_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_2_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_2_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed;
  reg        [2:0]    Lsu2Plugin_logic_lq_regs_2_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_2;
  wire                when_Lsu2Plugin_l338_2;
  reg                 Lsu2Plugin_logic_lq_regs_3_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_3_valid;
  reg                 Lsu2Plugin_logic_lq_regs_3_redo;
  reg                 Lsu2Plugin_logic_lq_regs_3_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_3_delete;
  reg                 Lsu2Plugin_logic_lq_regs_3_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_3_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_3_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_3_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed;
  reg        [2:0]    Lsu2Plugin_logic_lq_regs_3_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_3;
  wire                when_Lsu2Plugin_l338_3;
  reg                 Lsu2Plugin_logic_lq_regs_4_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_4_valid;
  reg                 Lsu2Plugin_logic_lq_regs_4_redo;
  reg                 Lsu2Plugin_logic_lq_regs_4_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_4_delete;
  reg                 Lsu2Plugin_logic_lq_regs_4_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_4_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_4_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_4_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed;
  reg        [2:0]    Lsu2Plugin_logic_lq_regs_4_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_4;
  wire                when_Lsu2Plugin_l338_4;
  reg                 Lsu2Plugin_logic_lq_regs_5_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_5_valid;
  reg                 Lsu2Plugin_logic_lq_regs_5_redo;
  reg                 Lsu2Plugin_logic_lq_regs_5_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_5_delete;
  reg                 Lsu2Plugin_logic_lq_regs_5_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_5_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_5_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_5_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed;
  reg        [2:0]    Lsu2Plugin_logic_lq_regs_5_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_5;
  wire                when_Lsu2Plugin_l338_5;
  reg                 Lsu2Plugin_logic_lq_regs_6_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_6_valid;
  reg                 Lsu2Plugin_logic_lq_regs_6_redo;
  reg                 Lsu2Plugin_logic_lq_regs_6_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_6_delete;
  reg                 Lsu2Plugin_logic_lq_regs_6_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_6_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_6_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_6_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed;
  reg        [2:0]    Lsu2Plugin_logic_lq_regs_6_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_6;
  wire                when_Lsu2Plugin_l338_6;
  reg                 Lsu2Plugin_logic_lq_regs_7_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_7_valid;
  reg                 Lsu2Plugin_logic_lq_regs_7_redo;
  reg                 Lsu2Plugin_logic_lq_regs_7_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_7_delete;
  reg                 Lsu2Plugin_logic_lq_regs_7_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_7_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_7_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_7_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed;
  reg        [2:0]    Lsu2Plugin_logic_lq_regs_7_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_7;
  wire                when_Lsu2Plugin_l338_7;
  reg        [6:0]    Lsu2Plugin_logic_lq_ptr_priority;
  reg        [6:0]    Lsu2Plugin_logic_lq_ptr_priorityLast;
  reg        [3:0]    Lsu2Plugin_logic_lq_ptr_alloc;
  reg        [3:0]    Lsu2Plugin_logic_lq_ptr_free;
  wire       [2:0]    Lsu2Plugin_logic_lq_ptr_allocReal;
  wire       [2:0]    Lsu2Plugin_logic_lq_ptr_freeReal;
  reg        [3:0]    Lsu2Plugin_logic_lq_tracker_freeNext;
  reg        [3:0]    Lsu2Plugin_logic_lq_tracker_free;
  reg        [0:0]    _zz_Lsu2Plugin_logic_lq_tracker_freeReduced;
  wire                when_UInt_l120;
  reg        [0:0]    Lsu2Plugin_logic_lq_tracker_freeReduced;
  wire       [0:0]    Lsu2Plugin_logic_lq_tracker_add;
  reg        [0:0]    Lsu2Plugin_logic_lq_tracker_sub;
  reg                 Lsu2Plugin_logic_lq_tracker_clear;
  wire                Lsu2Plugin_logic_lq_onCommit_lqAlloc_0;
  wire                Lsu2Plugin_logic_lq_onCommit_lqCommits_0;
  wire       [0:0]    Lsu2Plugin_logic_lq_onCommit_lqCommitCount;
  wire       [3:0]    Lsu2Plugin_logic_lq_onCommit_free;
  wire       [6:0]    Lsu2Plugin_logic_lq_onCommit_priority;
  wire                when_Lsu2Plugin_l454;
  wire                when_Lsu2Plugin_l454_1;
  wire                when_Lsu2Plugin_l454_2;
  wire                when_Lsu2Plugin_l454_3;
  wire                when_Lsu2Plugin_l454_4;
  wire                when_Lsu2Plugin_l454_5;
  wire                when_Lsu2Plugin_l454_6;
  wire                when_Lsu2Plugin_l454_7;
  reg                 Lsu2Plugin_logic_lq_reservation_kill;
  reg                 Lsu2Plugin_logic_lq_reservation_valid;
  reg        [31:0]   Lsu2Plugin_logic_lq_reservation_address;
  reg        [6:0]    Lsu2Plugin_logic_lq_reservation_counter;
  wire                when_Lsu2Plugin_l484;
  wire                Lsu2Plugin_logic_lq_hazardPrediction_hazard;
  reg                 Lsu2Plugin_logic_lq_hazardPrediction_write_valid;
  reg        [6:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address;
  reg        [2:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score;
  reg        [15:0]   Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag;
  reg        [2:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta;
  wire                Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_valid;
  wire       [6:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_address;
  wire       [2:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_score;
  wire       [15:0]   Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_tag;
  wire       [2:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_delta;
  wire                Lsu2Plugin_logic_lq_hitPrediction_hazard;
  wire                Lsu2Plugin_logic_lq_hitPrediction_write_valid;
  wire       [5:0]    Lsu2Plugin_logic_lq_hitPrediction_write_payload_address;
  wire       [5:0]    Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter;
  wire                Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_valid;
  wire       [5:0]    Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_address;
  wire       [5:0]    Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_data_counter;
  reg                 Lsu2Plugin_logic_sq_regs_0_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_0_valid;
  reg                 Lsu2Plugin_logic_sq_regs_0_redo;
  reg                 Lsu2Plugin_logic_sq_regs_0_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_0_delete;
  reg                 Lsu2Plugin_logic_sq_regs_0_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_0_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_0_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_0_commited;
  reg                 Lsu2Plugin_logic_sq_regs_0_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369;
  wire                when_Lsu2Plugin_l385;
  reg                 Lsu2Plugin_logic_sq_regs_1_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_1_valid;
  reg                 Lsu2Plugin_logic_sq_regs_1_redo;
  reg                 Lsu2Plugin_logic_sq_regs_1_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_1_delete;
  reg                 Lsu2Plugin_logic_sq_regs_1_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_1_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_1_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_1_commited;
  reg                 Lsu2Plugin_logic_sq_regs_1_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_1;
  wire                when_Lsu2Plugin_l385_1;
  reg                 Lsu2Plugin_logic_sq_regs_2_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_2_valid;
  reg                 Lsu2Plugin_logic_sq_regs_2_redo;
  reg                 Lsu2Plugin_logic_sq_regs_2_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_2_delete;
  reg                 Lsu2Plugin_logic_sq_regs_2_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_2_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_2_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_2_commited;
  reg                 Lsu2Plugin_logic_sq_regs_2_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_2;
  wire                when_Lsu2Plugin_l385_2;
  reg                 Lsu2Plugin_logic_sq_regs_3_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_3_valid;
  reg                 Lsu2Plugin_logic_sq_regs_3_redo;
  reg                 Lsu2Plugin_logic_sq_regs_3_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_3_delete;
  reg                 Lsu2Plugin_logic_sq_regs_3_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_3_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_3_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_3_commited;
  reg                 Lsu2Plugin_logic_sq_regs_3_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_3;
  wire                when_Lsu2Plugin_l385_3;
  reg                 Lsu2Plugin_logic_sq_regs_4_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_4_valid;
  reg                 Lsu2Plugin_logic_sq_regs_4_redo;
  reg                 Lsu2Plugin_logic_sq_regs_4_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_4_delete;
  reg                 Lsu2Plugin_logic_sq_regs_4_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_4_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_4_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_4_commited;
  reg                 Lsu2Plugin_logic_sq_regs_4_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_4;
  wire                when_Lsu2Plugin_l385_4;
  reg                 Lsu2Plugin_logic_sq_regs_5_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_5_valid;
  reg                 Lsu2Plugin_logic_sq_regs_5_redo;
  reg                 Lsu2Plugin_logic_sq_regs_5_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_5_delete;
  reg                 Lsu2Plugin_logic_sq_regs_5_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_5_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_5_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_5_commited;
  reg                 Lsu2Plugin_logic_sq_regs_5_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_5;
  wire                when_Lsu2Plugin_l385_5;
  reg                 Lsu2Plugin_logic_sq_regs_6_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_6_valid;
  reg                 Lsu2Plugin_logic_sq_regs_6_redo;
  reg                 Lsu2Plugin_logic_sq_regs_6_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_6_delete;
  reg                 Lsu2Plugin_logic_sq_regs_6_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_6_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_6_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_6_commited;
  reg                 Lsu2Plugin_logic_sq_regs_6_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_6;
  wire                when_Lsu2Plugin_l385_6;
  reg                 Lsu2Plugin_logic_sq_regs_7_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_7_valid;
  reg                 Lsu2Plugin_logic_sq_regs_7_redo;
  reg                 Lsu2Plugin_logic_sq_regs_7_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_7_delete;
  reg                 Lsu2Plugin_logic_sq_regs_7_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_7_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_7_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_7_commited;
  reg                 Lsu2Plugin_logic_sq_regs_7_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_7;
  wire                when_Lsu2Plugin_l385_7;
  reg                 Lsu2Plugin_logic_sq_mem_swap;
  reg        [2:0]    Lsu2Plugin_logic_sq_mem_op;
  reg        [5:0]    Lsu2Plugin_logic_sq_mem_physRd;
  reg                 Lsu2Plugin_logic_sq_mem_writeRd;
  reg        [6:0]    Lsu2Plugin_logic_sq_ptr_priority;
  reg        [6:0]    Lsu2Plugin_logic_sq_ptr_priorityLast;
  reg        [3:0]    Lsu2Plugin_logic_sq_ptr_alloc;
  reg        [3:0]    Lsu2Plugin_logic_sq_ptr_commit;
  reg        [3:0]    Lsu2Plugin_logic_sq_ptr_writeBack;
  reg        [3:0]    Lsu2Plugin_logic_sq_ptr_free;
  wire       [2:0]    Lsu2Plugin_logic_sq_ptr_allocReal;
  wire       [2:0]    Lsu2Plugin_logic_sq_ptr_freeReal /* verilator public */ ;
  wire       [2:0]    Lsu2Plugin_logic_sq_ptr_writeBackReal;
  wire       [2:0]    Lsu2Plugin_logic_sq_ptr_commitReal;
  wire       [3:0]    Lsu2Plugin_logic_sq_ptr_commitNext;
  reg                 Lsu2Plugin_logic_sq_ptr_onFree_valid;
  wire       [2:0]    Lsu2Plugin_logic_sq_ptr_onFree_payload;
  reg                 Lsu2Plugin_logic_sq_ptr_onFreeLast_valid;
  reg        [2:0]    Lsu2Plugin_logic_sq_ptr_onFreeLast_payload;
  wire                when_Lsu2Plugin_l572;
  wire       [3:0]    Lsu2Plugin_logic_sq_tracker_freeNext;
  reg        [3:0]    Lsu2Plugin_logic_sq_tracker_free;
  reg        [0:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeReduced;
  wire                when_UInt_l120_1;
  reg        [0:0]    Lsu2Plugin_logic_sq_tracker_freeReduced;
  reg        [0:0]    Lsu2Plugin_logic_sq_tracker_add;
  reg        [0:0]    Lsu2Plugin_logic_sq_tracker_sub;
  wire                Lsu2Plugin_logic_sq_onCommit_sqAlloc_0;
  wire       [0:0]    Lsu2Plugin_logic_sq_onCommit_sqCommits_0;
  wire       [3:0]    Lsu2Plugin_logic_sq_onCommit_commitComb;
  wire                when_Lsu2Plugin_l591;
  wire       [7:0]    _zz_44;
  wire                Lsu2Plugin_logic_allocation_loads_requests_0;
  wire       [0:0]    Lsu2Plugin_logic_allocation_loads_requestsCount;
  wire                Lsu2Plugin_logic_allocation_loads_full;
  wire       [3:0]    Lsu2Plugin_logic_allocation_loads_alloc;
  wire                Lsu2Plugin_logic_allocation_stores_requests_0;
  wire       [0:0]    Lsu2Plugin_logic_allocation_stores_requestsCount;
  wire                Lsu2Plugin_logic_allocation_stores_full;
  wire       [3:0]    Lsu2Plugin_logic_allocation_stores_alloc;
  wire                FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l620;
  wire                FrontendPlugin_dispatch_isFireing /* verilator public */ ;
  wire                Lsu2Plugin_logic_aguPush_0_pushLq;
  wire                Lsu2Plugin_logic_aguPush_0_pushSq;
  reg        [3:0]    _zz_Lsu2Plugin_logic_aguPush_0_dataMask;
  wire       [3:0]    Lsu2Plugin_logic_aguPush_0_dataMask;
  wire       [2:0]    switch_Utils_l1423;
  wire                Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_valid;
  wire       [6:0]    Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_payload;
  wire       [2:0]    Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
  wire       [15:0]   Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_tag;
  wire       [2:0]    Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_delta;
  wire       [21:0]   _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
  wire       [15:0]   Lsu2Plugin_logic_aguPush_0_hazardPrediction_hash;
  wire                Lsu2Plugin_logic_aguPush_0_hazardPrediction_hit;
  wire                Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_valid;
  wire       [5:0]    Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_payload;
  wire       [5:0]    Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
  wire                Lsu2Plugin_logic_aguPush_0_hitPrediction_likelyToHit;
  wire                when_Lsu2Plugin_l733;
  wire       [2:0]    switch_Utils_l1423_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_valid;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_input;
  wire       [6:0]    Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_priorityBits;
  wire       [14:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask;
  wire       [14:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_14;
  reg        [14:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_2_to_3;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_3;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_4_to_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_9;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_10_to_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_13;
  wire       [14:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pLow;
  wire       [6:0]    Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pHigh;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_input;
  wire       [6:0]    Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_priorityBits;
  wire       [14:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask;
  wire       [14:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_14;
  reg        [14:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_2_to_3;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_3;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_4_to_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_9;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_10_to_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_13;
  wire       [14:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pLow;
  wire       [6:0]    Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pHigh;
  wire       [7:0]    Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_1;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_3;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_7;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_8;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_9;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_1;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_3;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_7;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_8;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_9;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s1_valid;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_cmp;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_valid;
  reg                 _zz_Lsu2Plugin_logic_sharedPip_stages_1_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_valid;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_wake;
  reg                 Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap;
  reg                 Lsu2Plugin_logic_sharedPip_speculateHitTrapRecovered;
  reg                 Lsu2Plugin_logic_sharedPip_speculativeHitPredictionGotReschedule;
  reg                 Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled;
  reg                 Lsu2Plugin_logic_sharedPip_feed_takeAgu;
  wire                when_Lsu2Plugin_l830;
  wire                when_Lsu2Plugin_l831;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l834;
  reg                 Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask;
  reg                 Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask;
  wire                when_Lsu2Plugin_l838;
  wire                when_Lsu2Plugin_l839;
  wire                when_Lsu2Plugin_l841;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842;
  wire                when_Lsu2Plugin_l843;
  wire                when_Lsu2Plugin_l845;
  wire                when_Lsu2Plugin_l849;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC;
  wire                when_Lsu2Plugin_l920;
  wire                when_Lsu2Plugin_l929;
  wire       [2:0]    switch_Utils_l1423_2;
  wire       [2:0]    switch_Utils_l1423_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_isFireing;
  reg        [3:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT;
  wire                when_Lsu2Plugin_l959;
  wire                Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_valid;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_payload_robId;
  wire                Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_valid;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_payload_physical;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_haltRequest_Lsu2Plugin_l990;
  wire                when_Lsu2Plugin_l997;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_loopback;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_youngerMask;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_olderMaskEmpty;
  reg        [7:0]    Lsu2Plugin_logic_sharedPip_checkSqMask_hits;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_olderHit;
  wire       [7:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits;
  wire       [6:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask;
  wire       [14:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_14;
  reg        [14:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_10_to_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh;
  wire       [6:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pLow;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pHigh;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_4;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_5;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_6;
  wire       [2:0]    Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_isFireing;
  wire                when_Lsu2Plugin_l1046;
  wire                when_Lsu2Plugin_l1052;
  wire                Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_addressMatch;
  wire                Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_fullMatch;
  wire                Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_translationFailure;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_data;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_checkLqHits_endId;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_checkLqHits_startMask;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_checkLqHits_endMask;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_loopback;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMaskEmpty;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_hit;
  wire                when_Lsu2Plugin_l1104;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_hit;
  wire                when_Lsu2Plugin_l1104_1;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_hit;
  wire                when_Lsu2Plugin_l1104_2;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_hit;
  wire                when_Lsu2Plugin_l1104_3;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_hit;
  wire                when_Lsu2Plugin_l1104_4;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_hit;
  wire                when_Lsu2Plugin_l1104_5;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_hit;
  wire                when_Lsu2Plugin_l1104_6;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_hit;
  wire                when_Lsu2Plugin_l1104_7;
  wire                Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerHit;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_input;
  wire       [6:0]    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_priorityBits;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask;
  wire       [14:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_14;
  reg        [14:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_10_to_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pLow;
  wire       [6:0]    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pHigh;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_4;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_5;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_6;
  wire       [2:0]    Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel;
  reg                 Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress;
  reg                 Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_0;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_1;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_2;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted;
  wire                when_Lsu2Plugin_l1158;
  wire                _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
  reg        [31:0]   _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
  reg        [31:0]   _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_4;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_isFireing;
  wire                Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_valid /* verilator public */ ;
  wire                Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_isLoad /* verilator public */ ;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_address /* verilator public */ ;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_readData /* verilator public */ ;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_robId /* verilator public */ ;
  wire       [2:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_lqId /* verilator public */ ;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_size /* verilator public */ ;
  wire                Lsu2Plugin_logic_sharedPip_cacheRsp_doIt;
  reg                 Lsu2Plugin_logic_sharedPip_cacheRsp_success;
  wire                when_Lsu2Plugin_l1203;
  wire                when_Lsu2Plugin_l1205;
  wire                when_Lsu2Plugin_l1207;
  wire                when_Lsu2Plugin_l1209;
  wire                when_Lsu2Plugin_l1211;
  wire                when_Lsu2Plugin_l1213;
  wire       [2:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC;
  reg                 Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_valid;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_payload_robId;
  reg                 Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_payload_physical;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_ctrl_lqMask;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_ctrl_sqMask;
  reg                 Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
  wire                Lsu2Plugin_logic_sharedPip_ctrl_doCompletion;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_isFireing;
  wire                when_Lsu2Plugin_l1313;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
  wire                when_Lsu2Plugin_l1314;
  wire                when_Lsu2Plugin_l1333;
  wire                when_Lsu2Plugin_l1335;
  wire                _zz_when_Lsu2Plugin_l1348;
  reg        [2:0]    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score;
  wire                when_Lsu2Plugin_l1348;
  wire                when_Lsu2Plugin_l1351;
  wire                when_Lsu2Plugin_l1374;
  wire       [5:0]    _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next;
  wire       [6:0]    Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next;
  reg        [5:0]    _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter;
  wire                when_SInt_l131;
  wire                when_SInt_l132;
  wire                when_SInt_l138;
  reg                 Lsu2Plugin_logic_writeback_generation;
  reg        [1:0]    Lsu2Plugin_logic_writeback_waitOn_refillSlot;
  reg                 Lsu2Plugin_logic_writeback_waitOn_refillSlotAny;
  wire                Lsu2Plugin_logic_writeback_waitOn_ready;
  reg        [1:0]    Lsu2Plugin_logic_writeback_waitOn_refillSlotSet;
  reg                 Lsu2Plugin_logic_writeback_waitOn_refillSlotAnySet;
  wire                Lsu2Plugin_logic_writeback_feed_holdPrefetch;
  wire                toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_valid;
  wire                toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready;
  wire       [31:0]   toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_payload;
  reg                 toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rValid;
  reg        [31:0]   toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rData;
  wire                when_Stream_l369_2;
  wire                _zz_toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready;
  wire                Lsu2Plugin_logic_writeback_feed_prediction_valid;
  wire       [31:0]   Lsu2Plugin_logic_writeback_feed_prediction_payload;
  wire                Lsu2Plugin_logic_writeback_feed_io;
  wire       [1:0]    Lsu2Plugin_logic_writeback_feed_size;
  reg        [31:0]   Lsu2Plugin_logic_writeback_feed_data;
  reg                 Lsu2Plugin_logic_writeback_feed_skip;
  wire                Lsu2Plugin_logic_writeback_feed_doit;
  reg                 Lsu2Plugin_logic_writeback_feed_fire;
  reg        [3:0]    _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_valid;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_fault;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlot;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_generationKo;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_flush;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_prefetch;
  wire       [31:0]   Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_address;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_io;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_valid;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_fault;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlot;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_generationKo;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_flush;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_prefetch;
  wire       [31:0]   Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_address;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_io;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_valid;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_fault;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlot;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_generationKo;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_flush;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_prefetch;
  wire       [31:0]   Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_address;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_io;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_valid;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_fault;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_redo;
  reg        [1:0]    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlot;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlotAny;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_generationKo;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_flush;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_prefetch;
  reg        [31:0]   Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_address;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_io;
  reg                 Lsu2Plugin_logic_writeback_rsp_whitebox_valid /* verilator public */ ;
  wire                when_Lsu2Plugin_l1488;
  wire                when_Lsu2Plugin_l1498;
  wire                when_Lsu2Plugin_l1509;
  wire                when_Lsu2Plugin_l1521;
  wire                when_Lsu2Plugin_l1524;
  wire                when_Lsu2Plugin_l1524_1;
  wire                when_Lsu2Plugin_l1524_2;
  wire                when_Lsu2Plugin_l1524_3;
  wire                when_Lsu2Plugin_l1524_4;
  wire                when_Lsu2Plugin_l1524_5;
  wire                when_Lsu2Plugin_l1524_6;
  wire                when_Lsu2Plugin_l1524_7;
  reg                 Lsu2Plugin_logic_flush_busy;
  reg                 Lsu2Plugin_logic_flush_doit;
  reg                 Lsu2Plugin_logic_flush_withFree;
  reg        [2:0]    Lsu2Plugin_logic_flush_cmdPtr;
  reg        [2:0]    Lsu2Plugin_logic_flush_rspPtr;
  wire                FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548;
  wire                when_Lsu2Plugin_l1553;
  wire                Lsu2Plugin_setup_cacheStore_cmd_fire;
  wire                when_Lsu2Plugin_l1561;
  wire                when_Lsu2Plugin_l1569;
  wire                Lsu2Plugin_logic_special_lqOnTop;
  wire                Lsu2Plugin_logic_special_sqOnTop;
  wire                Lsu2Plugin_logic_special_storeWriteBackUsable;
  wire                Lsu2Plugin_logic_special_storeSpecial;
  wire                Lsu2Plugin_logic_special_loadSpecial;
  wire                Lsu2Plugin_logic_special_storeHit;
  wire                Lsu2Plugin_logic_special_loadHit;
  wire                Lsu2Plugin_logic_special_hit;
  reg                 LsuPlugin_peripheralBus_rsp_valid_regNext;
  reg                 Lsu2Plugin_logic_special_fire;
  reg                 Lsu2Plugin_logic_special_enabled;
  reg                 Lsu2Plugin_logic_special_isStore;
  reg                 Lsu2Plugin_logic_special_isLoad;
  reg                 Lsu2Plugin_logic_special_cmdSent;
  wire                LsuPlugin_peripheralBus_cmd_fire;
  reg        [3:0]    Lsu2Plugin_logic_special_robId /* verilator public */ ;
  reg        [5:0]    Lsu2Plugin_logic_special_loadPhysRd;
  reg        [31:0]   Lsu2Plugin_logic_special_loadAddress;
  reg        [31:0]   Lsu2Plugin_logic_special_loadAddressVirt;
  reg        [1:0]    Lsu2Plugin_logic_special_loadSize;
  reg                 Lsu2Plugin_logic_special_loadUnsigned;
  reg                 Lsu2Plugin_logic_special_loadWriteRd;
  reg        [31:0]   Lsu2Plugin_logic_special_storeAddress;
  reg        [31:0]   Lsu2Plugin_logic_special_storeAddressVirt;
  reg        [1:0]    Lsu2Plugin_logic_special_storeSize;
  reg        [31:0]   Lsu2Plugin_logic_special_storeData;
  reg        [3:0]    Lsu2Plugin_logic_special_storeMask;
  reg                 Lsu2Plugin_logic_special_storeAmo;
  reg                 Lsu2Plugin_logic_special_storeSc;
  wire       [31:0]   Lsu2Plugin_logic_special_address;
  wire       [31:0]   Lsu2Plugin_logic_special_addressVirt;
  wire                Lsu2Plugin_logic_special_isIo;
  wire                Lsu2Plugin_logic_special_isAtomic;
  reg                 Lsu2Plugin_logic_special_wakeRob_valid;
  wire       [3:0]    Lsu2Plugin_logic_special_wakeRob_payload_robId;
  reg                 Lsu2Plugin_logic_special_wakeRf_valid;
  wire       [5:0]    Lsu2Plugin_logic_special_wakeRf_payload_physical;
  wire                Lsu2Plugin_logic_special_atomic_wantExit;
  reg                 Lsu2Plugin_logic_special_atomic_wantStart;
  wire                Lsu2Plugin_logic_special_atomic_wantKill;
  reg        [31:0]   Lsu2Plugin_logic_special_atomic_readed;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1;
  wire                Lsu2Plugin_logic_special_atomic_alu_compare;
  wire                Lsu2Plugin_logic_special_atomic_alu_unsigned;
  wire       [31:0]   Lsu2Plugin_logic_special_atomic_alu_addSub;
  wire                Lsu2Plugin_logic_special_atomic_alu_less;
  wire                Lsu2Plugin_logic_special_atomic_alu_selectRf;
  wire       [2:0]    switch_Misc_l241_1;
  reg        [31:0]   Lsu2Plugin_logic_special_atomic_alu_raw;
  wire       [31:0]   Lsu2Plugin_logic_special_atomic_alu_result /* verilator public */ ;
  reg        [31:0]   Lsu2Plugin_logic_special_atomic_result;
  wire                when_Lsu2Plugin_l1683;
  wire                when_Lsu2Plugin_l1698;
  reg                 Lsu2Plugin_logic_special_atomic_gotReservation;
  reg        [1:0]    Lsu2Plugin_logic_special_atomic_lockDelayCounter;
  reg                 Lsu2Plugin_logic_special_atomic_comp_wakeRf;
  reg                 Lsu2Plugin_logic_special_atomic_comp_rfWrite;
  reg                 Lsu2Plugin_logic_special_atomic_loadWhitebox_valid /* verilator public */ ;
  wire       [31:0]   Lsu2Plugin_logic_special_atomic_loadWhitebox_readData /* verilator public */ ;
  reg                 Lsu2Plugin_logic_special_atomic_storeWhitebox_valid /* verilator public */ ;
  wire                Lsu2Plugin_logic_special_atomic_storeWhitebox_isSc /* verilator public */ ;
  wire                Lsu2Plugin_logic_special_atomic_storeWhitebox_scPassed /* verilator public */ ;
  wire                FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l1838;
  reg                 Lsu2Plugin_logic_lqFlush /* verilator public */ ;
  wire                when_Lsu2Plugin_l1913;
  wire                when_Lsu2Plugin_l1913_1;
  wire                when_Lsu2Plugin_l1913_2;
  wire                when_Lsu2Plugin_l1913_3;
  wire                when_Lsu2Plugin_l1913_4;
  wire                when_Lsu2Plugin_l1913_5;
  wire                when_Lsu2Plugin_l1913_6;
  wire                when_Lsu2Plugin_l1913_7;
  wire                sqAlloc_0_valid /* verilator public */ ;
  wire       [2:0]    sqAlloc_0_id /* verilator public */ ;
  wire                sqFree_valid /* verilator public */ ;
  wire       [2:0]    sqFree_payload /* verilator public */ ;
  wire       [32:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
  wire                EU0_BranchPlugin_logic_branch_badEarlyTaken;
  wire                EU0_ExecutionUnitBase_pipeline_execute_1_isFireing;
  wire                EU0_BranchPlugin_logic_branch_finalBranch_valid;
  wire       [1:0]    EU0_BranchPlugin_logic_branch_finalBranch_payload_address;
  wire       [31:0]   EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice;
  wire       [31:0]   EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget;
  wire                EU0_BranchPlugin_logic_branch_finalBranch_payload_data_taken;
  reg        [0:0]    MmuPlugin_logic_satp_mode;
  reg        [19:0]   MmuPlugin_logic_satp_ppn;
  reg                 MmuPlugin_logic_status_mxr;
  reg                 MmuPlugin_logic_status_sum;
  reg                 MmuPlugin_logic_status_mprv;
  wire       [0:0]    MmuPlugin_logic_satpModeWrite;
  reg                 FetchCachePlugin_setup_translationStorage_logic_refillOngoing;
  reg        [3:0]    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask;
  reg        [1:0]    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault;
  reg        [17:0]   FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willClear;
  reg        [1:0]    FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [1:0]    FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [1:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask;
  reg        [1:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault;
  reg        [7:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [9:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willClear;
  reg        [0:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_valueNext;
  reg        [0:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflow;
  reg                 Lsu2Plugin_setup_translationStorage_logic_refillOngoing;
  reg        [3:0]    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask;
  reg        [1:0]    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault;
  reg        [17:0]   Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willClear;
  reg        [1:0]    Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [1:0]    Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [1:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask;
  reg        [1:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault;
  reg        [7:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [9:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willClear;
  reg        [0:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_valueNext;
  reg        [0:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflow;
  reg                 Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg;
  wire                when_MmuPlugin_l278;
  reg                 Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg;
  wire                when_MmuPlugin_l278_1;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress;
  wire       [44:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid;
  wire       [44:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid;
  wire       [44:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid;
  wire       [44:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_translationPort_logic_read_1_readAddress;
  wire       [24:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid;
  wire       [24:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hit;
  wire       [5:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_4;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_5;
  reg        [5:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_1;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_2;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_3;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault;
  reg                 Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_needRefill;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_askRefill;
  wire                when_MmuPlugin_l315;
  wire                when_MmuPlugin_l316;
  wire                when_MmuPlugin_l318;
  wire                EU0_CsrAccessPlugin_logic_fsm_wantExit;
  reg                 EU0_CsrAccessPlugin_logic_fsm_wantStart;
  wire                EU0_CsrAccessPlugin_logic_fsm_wantKill;
  reg                 REG_CSR_773;
  reg                 REG_CSR_835;
  reg                 REG_CSR_833;
  reg                 REG_CSR_832;
  reg                 REG_CSR_3857;
  reg                 REG_CSR_3858;
  reg                 REG_CSR_3859;
  reg                 REG_CSR_3860;
  reg                 REG_CSR_769;
  reg                 REG_CSR_834;
  reg                 REG_CSR_768;
  reg                 REG_CSR_836;
  reg                 REG_CSR_772;
  reg                 REG_CSR_770;
  reg                 REG_CSR_771;
  reg                 REG_CSR_261;
  reg                 REG_CSR_323;
  reg                 REG_CSR_321;
  reg                 REG_CSR_320;
  reg                 REG_CSR_322;
  reg                 REG_CSR_256;
  reg                 REG_CSR_260;
  reg                 REG_CSR_324;
  reg                 REG_CSR_384;
  wire                CsrRamPlugin_setup_initPort_valid;
  wire                CsrRamPlugin_setup_initPort_ready;
  wire       [2:0]    CsrRamPlugin_setup_initPort_address;
  wire       [31:0]   CsrRamPlugin_setup_initPort_data;
  reg                 PrivilegedPlugin_setup_ramRead_valid;
  wire                PrivilegedPlugin_setup_ramRead_ready;
  reg        [2:0]    PrivilegedPlugin_setup_ramRead_address;
  wire       [31:0]   PrivilegedPlugin_setup_ramRead_data;
  reg                 PrivilegedPlugin_setup_ramWrite_valid;
  wire                PrivilegedPlugin_setup_ramWrite_ready;
  reg        [2:0]    PrivilegedPlugin_setup_ramWrite_address;
  reg        [31:0]   PrivilegedPlugin_setup_ramWrite_data;
  wire                EU0_CsrAccessPlugin_logic_ramReadPort_valid;
  wire                EU0_CsrAccessPlugin_logic_ramReadPort_ready;
  wire       [2:0]    EU0_CsrAccessPlugin_logic_ramReadPort_address;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_ramReadPort_data;
  wire                EU0_CsrAccessPlugin_logic_ramWritePort_valid;
  wire                EU0_CsrAccessPlugin_logic_ramWritePort_ready;
  wire       [2:0]    EU0_CsrAccessPlugin_logic_ramWritePort_address;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_ramWritePort_data;
  reg        [3:0]    CsrRamPlugin_logic_flush_counter;
  wire                CsrRamPlugin_logic_flush_done;
  wire                when_CsrRamPlugin_l61;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits;
  wire                CsrRamPlugin_logic_writeLogic_hit;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_input;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_oh;
  wire                _zz_PrivilegedPlugin_setup_ramWrite_ready;
  wire                _zz_CsrRamPlugin_setup_initPort_ready;
  wire       [1:0]    CsrRamPlugin_logic_writeLogic_sel;
  wire                CsrRamPlugin_logic_writeLogic_port_valid;
  wire       [2:0]    CsrRamPlugin_logic_writeLogic_port_payload_address;
  wire       [31:0]   CsrRamPlugin_logic_writeLogic_port_payload_data;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits;
  wire                CsrRamPlugin_logic_readLogic_hit;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_input;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_oh;
  wire                _zz_PrivilegedPlugin_setup_ramRead_ready;
  wire       [0:0]    CsrRamPlugin_logic_readLogic_sel;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_port_address;
  wire       [31:0]   CsrRamPlugin_logic_readLogic_port_data;
  reg                 PrivilegedPlugin_logic_interrupt_valid;
  reg        [3:0]    PrivilegedPlugin_logic_interrupt_code;
  reg        [1:0]    PrivilegedPlugin_logic_interrupt_targetPrivilege;
  wire                when_PrivilegedPlugin_l638;
  wire                when_PrivilegedPlugin_l638_1;
  wire                when_PrivilegedPlugin_l644;
  wire                when_PrivilegedPlugin_l644_1;
  wire                when_PrivilegedPlugin_l644_2;
  wire                when_PrivilegedPlugin_l644_3;
  wire                when_PrivilegedPlugin_l644_4;
  wire                when_PrivilegedPlugin_l644_5;
  wire                when_PrivilegedPlugin_l644_6;
  wire                when_PrivilegedPlugin_l644_7;
  wire                when_PrivilegedPlugin_l644_8;
  reg                 PrivilegedPlugin_logic_decoderInterrupt_raised;
  reg                 PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt;
  reg        [2:0]    PrivilegedPlugin_logic_decoderInterrupt_counter;
  wire                PrivilegedPlugin_logic_decoderInterrupt_doIt;
  wire                when_PrivilegedPlugin_l675;
  wire                when_PrivilegedPlugin_l679;
  wire                PrivilegedPlugin_logic_decoderInterrupt_buffer_sample;
  reg        [3:0]    PrivilegedPlugin_logic_decoderInterrupt_buffer_code;
  reg        [1:0]    PrivilegedPlugin_logic_decoderInterrupt_buffer_targetPrivilege;
  reg        [1:0]    PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped;
  reg        [3:0]    PrivilegedPlugin_logic_exception_code;
  wire                when_PrivilegedPlugin_l696;
  wire                when_PrivilegedPlugin_l709;
  wire                when_PrivilegedPlugin_l709_1;
  wire                when_PrivilegedPlugin_l709_2;
  wire                when_PrivilegedPlugin_l709_3;
  wire                when_PrivilegedPlugin_l709_4;
  wire                when_PrivilegedPlugin_l709_5;
  wire                when_PrivilegedPlugin_l709_6;
  wire       [1:0]    PrivilegedPlugin_logic_exception_targetPrivilege;
  wire                PrivilegedPlugin_logic_fsm_wantExit;
  reg                 PrivilegedPlugin_logic_fsm_wantStart;
  wire                PrivilegedPlugin_logic_fsm_wantKill;
  reg                 PrivilegedPlugin_logic_fsm_trap_fire;
  reg                 PrivilegedPlugin_logic_fsm_trap_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_fsm_trap_code;
  reg        [1:0]    PrivilegedPlugin_logic_fsm_trap_targetPrivilege;
  wire       [1:0]    PrivilegedPlugin_logic_fsm_xret_sourcePrivilege;
  reg        [1:0]    PrivilegedPlugin_logic_fsm_xret_targetPrivilege;
  wire                FetchPlugin_stages_0_haltRequest_PrivilegedPlugin_l975;
  wire                trap_fire /* verilator public */ ;
  wire       [3:0]    trap_code /* verilator public */ ;
  wire                trap_interrupt /* verilator public */ ;
  wire       [31:0]   trap_tval /* verilator public */ ;
  reg        [2:0]    EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_ramSel;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_regs_microOp;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_doImm;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_doMask;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_doClear;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_regs_rs1;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_implemented;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_trap;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_flushPipeline;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_read;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_write;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_regs_aluInput;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_regs_csrValue;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_immZero;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_srcZero;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_csrWrite;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_csrRead;
  wire                COMB_CSR_773;
  wire                COMB_CSR_835;
  wire                COMB_CSR_833;
  wire                COMB_CSR_832;
  wire                COMB_CSR_3857;
  wire                COMB_CSR_3858;
  wire                COMB_CSR_3859;
  wire                COMB_CSR_3860;
  wire                COMB_CSR_769;
  wire                COMB_CSR_834;
  wire                COMB_CSR_768;
  wire                COMB_CSR_836;
  wire                COMB_CSR_772;
  wire                COMB_CSR_770;
  wire                COMB_CSR_771;
  wire                COMB_CSR_261;
  wire                COMB_CSR_323;
  wire                COMB_CSR_321;
  wire                COMB_CSR_320;
  wire                COMB_CSR_322;
  wire                COMB_CSR_256;
  wire                COMB_CSR_260;
  wire                COMB_CSR_324;
  wire                COMB_CSR_384;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_trap;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_write;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_read;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_onDecodeDo;
  wire                when_CsrAccessPlugin_l183;
  wire                when_MmuPlugin_l218;
  reg                 EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  reg                 EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire                when_CsrAccessPlugin_l272;
  wire                when_CsrAccessPlugin_l278;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_masked;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
  reg                 EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  reg                 EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo;
  wire                when_CsrAccessPlugin_l327;
  wire                when_CsrAccessPlugin_l328;
  wire                when_CsrAccessPlugin_l328_1;
  wire                when_CsrAccessPlugin_l328_2;
  wire                when_CsrAccessPlugin_l328_3;
  wire                when_CsrAccessPlugin_l328_4;
  wire                when_CsrAccessPlugin_l328_5;
  wire                when_CsrAccessPlugin_l327_1;
  wire                when_CsrAccessPlugin_l328_6;
  wire                when_CsrAccessPlugin_l328_7;
  wire                when_CsrAccessPlugin_l328_8;
  wire                when_CsrAccessPlugin_l328_9;
  wire                when_CsrAccessPlugin_l333;
  wire                when_CsrAccessPlugin_l328_10;
  reg                 EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired;
  wire                when_CsrAccessPlugin_l338;
  wire                when_CsrAccessPlugin_l342;
  reg                 EU0_CsrAccessPlugin_logic_fsm_isDone;
  reg                 EU0_CsrAccessPlugin_logic_fsm_isCompletionReady;
  reg        [2:0]    EU0_CsrAccessPlugin_logic_fsm_stateReg;
  reg        [2:0]    EU0_CsrAccessPlugin_logic_fsm_stateNext;
  wire       [11:0]   switch_CsrAccessPlugin_l206;
  wire                when_CsrAccessPlugin_l285;
  wire                when_CsrAccessPlugin_l311;
  wire                EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_CsrAccessPlugin_l375;
  wire                when_CsrAccessPlugin_l378;
  wire                csrAccess_valid /* verilator public */ ;
  wire       [3:0]    csrAccess_payload_robId /* verilator public */ ;
  wire       [11:0]   csrAccess_payload_address /* verilator public */ ;
  wire       [31:0]   csrAccess_payload_write /* verilator public */ ;
  wire       [31:0]   csrAccess_payload_read /* verilator public */ ;
  wire                csrAccess_payload_writeDone /* verilator public */ ;
  wire                csrAccess_payload_readDone /* verilator public */ ;
  wire                csrAccess_payload_fsDirty /* verilator public */ ;
  wire                EU0_ExecutionUnitBase_pipeline_execute_2_isFireing;
  wire       [1:0]    EnvCallPlugin_logic_xretPriv;
  reg                 EnvCallPlugin_logic_trap;
  wire                when_EnvCallPlugin_l99;
  wire                when_EnvCallPlugin_l100;
  wire                when_EnvCallPlugin_l108;
  wire                when_EnvCallPlugin_l112;
  wire                when_EnvCallPlugin_l113;
  wire                EnvCallPlugin_logic_flushes_wantExit;
  reg                 EnvCallPlugin_logic_flushes_wantStart;
  wire                EnvCallPlugin_logic_flushes_wantKill;
  wire                FetchPlugin_stages_0_haltRequest_EnvCallPlugin_l138;
  reg                 EnvCallPlugin_logic_flushes_vmaInv;
  reg                 EnvCallPlugin_logic_flushes_fetchInv;
  reg                 EnvCallPlugin_logic_flushes_flushData;
  reg        [2:0]    EnvCallPlugin_logic_flushes_stateReg;
  reg        [2:0]    EnvCallPlugin_logic_flushes_stateNext;
  wire                when_EnvCallPlugin_l148;
  wire                when_MmuPlugin_l356;
  reg                 FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg;
  wire                when_MmuPlugin_l278_2;
  wire       [1:0]    FetchCachePlugin_logic_translationPort_logic_read_0_readAddress;
  wire       [44:0]   _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid;
  wire       [44:0]   _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid;
  wire       [44:0]   _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid;
  wire       [44:0]   _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid;
  wire       [1:0]    FetchCachePlugin_logic_translationPort_logic_read_1_readAddress;
  wire       [24:0]   _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid;
  wire       [24:0]   _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid;
  wire       [5:0]    FetchCachePlugin_logic_translationPort_logic_ctrl_hits;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hit;
  wire       [5:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_4;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_5;
  reg        [5:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_1;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_2;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_3;
  wire       [5:0]    FetchCachePlugin_logic_translationPort_logic_ctrl_oh;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineException;
  wire       [31:0]   FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault;
  reg                 FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_needRefill;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_askRefill;
  wire                when_MmuPlugin_l315_1;
  wire                when_MmuPlugin_l316_1;
  wire                when_MmuPlugin_l356_1;
  wire                MmuPlugin_logic_refill_wantExit;
  reg                 MmuPlugin_logic_refill_wantStart;
  wire                MmuPlugin_logic_refill_wantKill;
  wire                MmuPlugin_logic_refill_busy;
  reg        [1:0]    MmuPlugin_logic_refill_portOhReg;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask;
  reg        [31:0]   MmuPlugin_logic_refill_virtual;
  wire       [1:0]    MmuPlugin_logic_refill_portsRequests;
  reg                 MmuPlugin_logic_refill_portsRequest;
  wire       [1:0]    MmuPlugin_logic_refill_portsRequests_ohFirst_input;
  wire       [1:0]    MmuPlugin_logic_refill_portsRequests_ohFirst_masked;
  wire       [1:0]    MmuPlugin_logic_refill_portsOh;
  reg        [1:0]    MmuPlugin_logic_refill_portsOh_regNext;
  reg        [31:0]   _zz_MmuPlugin_logic_refill_portsAddress;
  reg        [31:0]   _zz_MmuPlugin_logic_refill_portsAddress_1;
  wire       [31:0]   MmuPlugin_logic_refill_portsAddress;
  reg        [1:0]    MmuPlugin_logic_refill_cacheRefill;
  reg                 MmuPlugin_logic_refill_cacheRefillAny;
  reg        [1:0]    MmuPlugin_logic_refill_cacheRefillSet;
  reg                 MmuPlugin_logic_refill_cacheRefillAnySet;
  wire                MmuPlugin_logic_refill_doWake;
  reg        [31:0]   MmuPlugin_logic_refill_load_address;
  reg                 MmuPlugin_logic_refill_load_rsp_valid;
  reg        [31:0]   MmuPlugin_logic_refill_load_rsp_payload_data;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_fault;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_redo;
  reg        [1:0]    MmuPlugin_logic_refill_load_rsp_payload_refillSlot;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_refillSlotAny;
  wire       [31:0]   MmuPlugin_logic_refill_load_readed;
  wire                when_MmuPlugin_l418;
  wire                MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_flags_R;
  wire                MmuPlugin_logic_refill_load_flags_W;
  wire                MmuPlugin_logic_refill_load_flags_X;
  wire                MmuPlugin_logic_refill_load_flags_U;
  wire                MmuPlugin_logic_refill_load_flags_G;
  wire                MmuPlugin_logic_refill_load_flags_A;
  wire                MmuPlugin_logic_refill_load_flags_D;
  wire       [31:0]   _zz_MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_leaf;
  reg                 MmuPlugin_logic_refill_load_exception;
  reg        [31:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_0;
  reg        [31:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_1;
  wire                MmuPlugin_logic_refill_load_levelException_0;
  reg                 MmuPlugin_logic_refill_load_levelException_1;
  reg        [31:0]   MmuPlugin_logic_refill_load_nextLevelBase;
  wire                when_MmuPlugin_l446;
  reg                 MmuPlugin_logic_invalidate_requested;
  reg                 MmuPlugin_logic_invalidate_canStart;
  reg        [2:0]    MmuPlugin_logic_invalidate_counter;
  wire                MmuPlugin_logic_invalidate_done;
  wire                when_MmuPlugin_l522;
  wire                FetchPlugin_stages_0_haltRequest_MmuPlugin_l533;
  wire                when_MmuPlugin_l535;
  wire                when_MmuPlugin_l541;
  reg                 MmuPlugin_logic_invalidate_done_regNext;
  wire                when_MmuPlugin_l545;
  wire                when_Pipeline_l278;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s0_ready_output;
  wire                when_Pipeline_l278_1;
  wire                when_Connection_l74;
  reg        [9:0]    Lsu2Plugin_logic_special_atomic_stateReg;
  reg        [9:0]    Lsu2Plugin_logic_special_atomic_stateNext;
  wire                when_Lsu2Plugin_l1704;
  wire                when_Lsu2Plugin_l1705;
  wire                Lsu2Plugin_setup_cacheLoad_cmd_fire;
  wire                when_Lsu2Plugin_l1715;
  wire                when_Lsu2Plugin_l1828;
  wire                when_StateMachine_l253;
  wire                when_StateMachine_l253_1;
  reg        [2:0]    MmuPlugin_logic_refill_stateReg;
  reg        [2:0]    MmuPlugin_logic_refill_stateNext;
  wire                when_MmuPlugin_l482;
  wire                when_MmuPlugin_l482_1;
  wire                when_MmuPlugin_l491;
  wire                when_MmuPlugin_l499;
  wire                DecoderPlugin_logic_slots_0_rdZero;
  wire                _zz_FrontendPlugin_decoded_SQ_ALLOC_0;
  wire                _zz_FrontendPlugin_decoded_SQ_ALLOC_0_1;
  reg                 DecoderPlugin_logic_slots_0_x0AlwaysZero;
  wire                _zz_FrontendPlugin_decoded_WRITE_RD_0;
  wire                DecoderPlugin_logic_exception_set;
  wire                DecoderPlugin_logic_exception_clear;
  reg                 DecoderPlugin_logic_exception_trigged;
  wire                when_DecoderPlugin_l302;
  reg                 DecoderPlugin_logic_exception_exceptionReg_0;
  wire                when_DecoderPlugin_l303;
  reg                 DecoderPlugin_logic_exception_fetchFaultReg_0;
  wire                when_DecoderPlugin_l304;
  reg                 DecoderPlugin_logic_exception_fetchFaultPageReg_0;
  wire                when_DecoderPlugin_l306;
  reg                 DecoderPlugin_logic_exception_debugEnterReg_0;
  wire                when_DecoderPlugin_l307;
  reg        [31:0]   DecoderPlugin_logic_exception_epcReg_0;
  wire                when_DecoderPlugin_l308;
  reg        [31:0]   DecoderPlugin_logic_exception_instReg_0;
  wire                when_DecoderPlugin_l309;
  reg                 DecoderPlugin_logic_exception_compressedFaultReg_0;
  wire                DecoderPlugin_logic_exception_compressedFault;
  wire                DecoderPlugin_logic_exception_fetchFault;
  wire                DecoderPlugin_logic_exception_fetchFaultPage;
  wire                DecoderPlugin_logic_exception_debugEnter;
  wire       [31:0]   DecoderPlugin_logic_exception_pc;
  wire                DecoderPlugin_logic_exception_pipelineEmpty;
  wire                DecoderPlugin_logic_exception_doIt;
  reg                 DecoderPlugin_logic_exception_doItAgain;
  wire                _zz_FrontendPlugin_decoded_isFlushingRoot;
  wire                FrontendPlugin_decoded_haltRequest_DecoderPlugin_l324;
  wire                FrontendPlugin_decoded_haltRequest_DecoderPlugin_l325;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_1;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_2;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_3;
  wire                switch_Misc_l241_2;
  reg        [31:0]   _zz_FrontendPlugin_decoded_OFFSET_0;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rs1Link;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdEquRs1;
  wire       [1:0]    DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_0_applyIt_badTaken;
  wire                when_DecoderPredictionPlugin_l212;
  wire                when_DecoderPredictionPlugin_l213;
  wire                when_DecoderPredictionPlugin_l219;
  wire                DecoderPredictionPlugin_logic_decodePatch_applyIt_hit;
  wire                FrontendPlugin_serialized_isFireing;
  reg                 DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle;
  wire                when_DecoderPredictionPlugin_l236;
  wire                when_DecoderPredictionPlugin_l243;
  wire                when_DecoderPredictionPlugin_l244;
  wire                ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                ALU0_ExecutionUnitBase_pipeline_push_port_valid;
  wire       [3:0]    ALU0_ExecutionUnitBase_pipeline_push_port_robId;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_push_port_physRd;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2;
  wire                ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  wire       [3:0]    ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  wire                ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid;
  wire       [3:0]    ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_isFireing;
  wire                EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                EU0_ExecutionUnitBase_pipeline_push_port_valid;
  wire                EU0_ExecutionUnitBase_pipeline_push_port_ready;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_push_port_robId;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_push_port_physRd;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_push_port_context_0;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_push_port_context_1;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD;
  wire                EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid;
  wire                EU0_ExecutionUnitBase_pipeline_writeBack_0_write_ready;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  wire                EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_ExecutionUnitBase_l303;
  wire                EU0_ExecutionUnitBase_pipeline_completion_0_port_valid;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  wire                EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_fire;
  wire                EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_valid;
  wire       [3:0]    EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_payload_robId;
  wire                EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_fire;
  wire                EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_valid;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_payload_physical;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_ready_output;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_0_ready_output;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_1_ready_output;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_1_ready;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output;
  wire                when_Pipeline_l278_2;
  wire                when_Pipeline_l278_3;
  wire                when_Pipeline_l278_4;
  wire                when_Connection_l74_1;
  wire                when_Connection_l74_2;
  wire                when_Connection_l74_3;
  wire                BranchContextPlugin_free_dispatchMem_writes_0_port_valid;
  wire       [1:0]    BranchContextPlugin_free_dispatchMem_writes_0_port_payload_address;
  wire       [26:0]   BranchContextPlugin_free_dispatchMem_writes_0_port_payload_data;
  wire                BranchContextPlugin_free_learn_valid;
  wire       [1:0]    BranchContextPlugin_free_learn_bid;
  wire       [64:0]   _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice;
  wire       [26:0]   BranchContextPlugin_free_learn_raw;
  wire       [7:0]    DispatchPlugin_logic_queueStaticWakeTransposed_0;
  wire       [7:0]    DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0;
  reg        [3:0]    DispatchPlugin_logic_ptr_next;
  reg        [3:0]    DispatchPlugin_logic_ptr_current;
  wire                toplevel_DispatchPlugin_logic_queue_io_push_fire;
  wire                FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l187;
  wire                DispatchPlugin_logic_push_skip;
  wire                DispatchPlugin_logic_push_fenceOlder;
  wire                DispatchPlugin_logic_push_fenceYounger;
  wire                when_DispatchPlugin_l192;
  reg                 DispatchPlugin_logic_push_fenceYoungerLast;
  wire                DispatchPlugin_logic_push_commitNotWaitingOnUs;
  wire                FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l195;
  wire                FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l196;
  wire       [7:0]    DispatchPlugin_logic_push_slots_0_self;
  wire       [7:0]    DispatchPlugin_logic_push_slots_0_events_0;
  wire       [7:0]    DispatchPlugin_logic_push_slots_0_events_1;
  wire                DispatchPlugin_logic_pop_0_stagesList_0_valid;
  reg                 DispatchPlugin_logic_pop_0_stagesList_1_valid;
  wire       [7:0]    DispatchPlugin_logic_pop_0_portEventFull;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_1;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_2;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_4;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_5;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_6;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3;
  wire                toplevel_DispatchPlugin_logic_queue_io_schedules_0_fire;
  wire       [7:0]    DispatchPlugin_logic_pop_0_wake_L0_mask;
  wire                DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid;
  wire       [5:0]    DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical;
  wire                DispatchPlugin_logic_pop_1_stagesList_0_valid;
  reg                 DispatchPlugin_logic_pop_1_stagesList_1_valid;
  wire       [7:0]    DispatchPlugin_logic_pop_1_portEventFull;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_1;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_2;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_4;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_5;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_6;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_0;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_1;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_2;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_3;
  wire                DispatchPlugin_logic_pop_1_stagesList_1_haltRequest_DispatchPlugin_l292;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_0;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_1;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_2;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_3;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_0;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_1;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_2;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_3;
  reg                 DispatchPlugin_logic_pop_1_stagesList_0_ready_output;
  wire                when_Pipeline_l278_5;
  wire                when_Connection_l74_4;
  wire                DispatchPlugin_logic_wake_dynamic_offseted_0_valid;
  wire       [2:0]    DispatchPlugin_logic_wake_dynamic_offseted_0_payload;
  wire                DispatchPlugin_logic_wake_dynamic_offseted_1_valid;
  wire       [2:0]    DispatchPlugin_logic_wake_dynamic_offseted_1_payload;
  wire                DispatchPlugin_logic_wake_dynamic_offseted_2_valid;
  wire       [2:0]    DispatchPlugin_logic_wake_dynamic_offseted_2_payload;
  wire                DispatchPlugin_logic_wake_dynamic_offseted_3_valid;
  wire       [2:0]    DispatchPlugin_logic_wake_dynamic_offseted_3_payload;
  wire       [7:0]    DispatchPlugin_logic_wake_dynamic_masks_0;
  wire       [7:0]    DispatchPlugin_logic_wake_dynamic_masks_1;
  wire       [7:0]    DispatchPlugin_logic_wake_dynamic_masks_2;
  wire       [7:0]    DispatchPlugin_logic_wake_dynamic_masks_3;
  wire       [7:0]    DispatchPlugin_logic_wake_statics_0_popMask;
  wire       [7:0]    DispatchPlugin_logic_wake_statics_0_history_0;
  (* keep , syn_keep *) wire       [7:0]    DispatchPlugin_logic_wake_optReduce_relaxed /* synthesis syn_keep = 1 */ ;
  wire       [7:0]    DispatchPlugin_logic_wake_optReduce_reduced;
  wire                DispatchPlugin_logic_whitebox_issuePorts_0_valid /* verilator public */ ;
  wire       [3:0]    DispatchPlugin_logic_whitebox_issuePorts_0_payload_robId /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_0_payload_physRd /* verilator public */ ;
  wire                DispatchPlugin_logic_whitebox_issuePorts_1_valid /* verilator public */ ;
  wire       [3:0]    DispatchPlugin_logic_whitebox_issuePorts_1_payload_robId /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_1_payload_physRd /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_1_payload_context_0 /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_1_payload_context_1 /* verilator public */ ;
  wire                integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  wire       [3:0]    integer_RegFilePlugin_logic_writeMerges_0_bus_robId;
  wire       [1:0]    _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0;
  wire                _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_1;
  reg        [1:0]    _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_2;
  wire                integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0;
  wire                integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_1;
  wire       [1:0]    _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_3;
  wire                integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data;
  wire                integer_RegFilePlugin_logic_writeMerges_1_bus_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_1_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_1_bus_data;
  wire       [3:0]    integer_RegFilePlugin_logic_writeMerges_1_bus_robId;
  wire                integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                when_RegFilePlugin_l327;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                when_RegFilePlugin_l327_1;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                when_RegFilePlugin_l327_2;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                when_RegFilePlugin_l327_3;
  wire                integer_write_0_valid /* verilator public */ ;
  wire       [5:0]    integer_write_0_address /* verilator public */ ;
  wire       [31:0]   integer_write_0_data /* verilator public */ ;
  wire       [3:0]    integer_write_0_robId /* verilator public */ ;
  wire                integer_write_1_valid /* verilator public */ ;
  wire       [5:0]    integer_write_1_address /* verilator public */ ;
  wire       [31:0]   integer_write_1_data /* verilator public */ ;
  wire       [3:0]    integer_write_1_robId /* verilator public */ ;
  wire                RobPlugin_logic_completionMem_targetWrite_valid;
  wire       [3:0]    RobPlugin_logic_completionMem_targetWrite_payload_address;
  wire       [0:0]    RobPlugin_logic_completionMem_targetWrite_payload_data;
  wire       [3:0]    RobPlugin_logic_completionMem_init_0_robId;
  wire       [3:0]    RobPlugin_logic_completionMem_reads_0_targetRead_address;
  wire       [0:0]    RobPlugin_logic_completionMem_reads_0_targetRead_data;
  wire       [3:0]    _zz_CommitPlugin_setup_robLineMask_mask;
  wire       [3:0]    _zz_when_RobPlugin_l118;
  wire                when_RobPlugin_l118;
  wire                when_RobPlugin_l118_1;
  wire                when_RobPlugin_l118_2;
  wire                when_RobPlugin_l118_3;
  wire                when_RobPlugin_l123;
  wire       [3:0]    _zz_CommitPlugin_logic_commit_active;
  wire       [3:0]    _zz_integer_RfAllocationPlugin_logic_push_mask_0;
  wire       [3:0]    _zz_commit_pc_0;
  wire       [3:0]    _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire       [3:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0;
  wire       [3:0]    _zz_integer_RfAllocationPlugin_logic_push_writeRd_0;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire       [3:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0;
  wire       [3:0]    _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0;
  wire       [3:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0;
  wire       [3:0]    _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0;
  wire       [3:0]    _zz_BranchContextPlugin_logic_onCommit_isBranch_0;
  wire       [3:0]    _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0;
  wire       [3:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch;
  wire       [3:0]    _zz_HistoryPlugin_logic_onCommit_isTaken_0;
  wire       [3:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken;
  wire       [3:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_healPush;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID;
  wire       [3:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB;
  wire                RobPlugin_logic_whitebox_completionsPorts_0_valid /* verilator public */ ;
  wire       [3:0]    RobPlugin_logic_whitebox_completionsPorts_0_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_1_valid /* verilator public */ ;
  wire       [3:0]    RobPlugin_logic_whitebox_completionsPorts_1_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_2_valid /* verilator public */ ;
  wire       [3:0]    RobPlugin_logic_whitebox_completionsPorts_2_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_3_valid /* verilator public */ ;
  wire       [3:0]    RobPlugin_logic_whitebox_completionsPorts_3_payload_id /* verilator public */ ;
  reg        [6:0]    RfDependencyPlugin_logic_forRf_integer_init_counter;
  wire                RfDependencyPlugin_logic_forRf_integer_init_busy;
  reg                 _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0;
  reg        [3:0]    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0;
  wire                when_RfDependencyPlugin_l228;
  wire                when_RfDependencyPlugin_l232;
  reg                 _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0;
  reg        [3:0]    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0;
  wire                when_RfDependencyPlugin_l228_1;
  wire                when_RfDependencyPlugin_l232_1;
  reg                 FrontendPlugin_allocated_ready_output;
  wire                FrontendPlugin_serialized_ready_output;
  wire                when_Connection_l66;
  reg                 FrontendPlugin_decoded_ready_output;
  wire                _zz_FrontendPlugin_decompressed_isFlushed;
  wire                FrontendPlugin_decompressed_ready_output;
  wire                FrontendPlugin_decompressed_ready;
  wire                FrontendPlugin_aligned_ready_output;
  wire                when_Pipeline_l278_6;
  wire                when_Pipeline_l278_7;
  wire                when_Pipeline_l278_8;
  wire                when_Connection_l74_5;
  wire                when_Connection_l74_6;
  reg        [6:0]    PcPlugin_logic_init_counter;
  wire                PcPlugin_logic_init_booted;
  wire                PcPlugin_logic_fetchPc_output_valid;
  wire                PcPlugin_logic_fetchPc_output_ready;
  wire       [31:0]   PcPlugin_logic_fetchPc_output_payload;
  reg        [31:0]   PcPlugin_logic_fetchPc_pcReg /* verilator public */ ;
  reg                 PcPlugin_logic_fetchPc_correction;
  reg                 PcPlugin_logic_fetchPc_correctionReg;
  wire                PcPlugin_logic_fetchPc_output_fire;
  wire                PcPlugin_logic_fetchPc_corrected;
  wire                PcPlugin_logic_fetchPc_pcRegPropagate;
  reg                 PcPlugin_logic_fetchPc_inc;
  wire                when_PcPlugin_l84;
  wire                when_PcPlugin_l84_1;
  reg        [31:0]   PcPlugin_logic_fetchPc_pc;
  reg                 PcPlugin_logic_fetchPc_flushed;
  wire                when_PcPlugin_l100;
  wire                PcPlugin_logic_fetchPc_fetcherHalt;
  wire                fetchLastFire /* verilator public */ ;
  wire       [11:0]   fetchLastId /* verilator public */ ;
  wire                FetchPlugin_stages_2_ready_output;
  wire                when_Connection_l66_1;
  reg                 FetchPlugin_stages_1_ready_output;
  wire                when_Connection_l54;
  reg                 FetchPlugin_stages_0_ready_output;
  wire                when_Pipeline_l278_9;
  wire                when_Pipeline_l278_10;
  wire                when_Connection_l74_7;
  wire                when_Connection_l74_8;
  reg                 FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_WORD_s2mBuffer;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_FETCH_PC_s2mBuffer;
  reg                 FetchPlugin_stages_2_Fetch_WORD_FAULT_s2mBuffer;
  reg                 FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE_s2mBuffer;
  reg        [23:0]   FetchPlugin_stages_2_BRANCH_HISTORY_s2mBuffer;
  reg        [11:0]   FetchPlugin_stages_2_FETCH_ID_s2mBuffer;
  reg                 FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID_s2mBuffer;
  reg        [0:0]    FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT_s2mBuffer;
  reg        [31:0]   FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT_s2mBuffer;
  reg                 FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID_s2mBuffer;
  reg                 FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE_s2mBuffer;
  reg        [1:0]    FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_0;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_FETCH_PC_INC_s2mBuffer;
  reg        [3:0]    PrivilegedPlugin_logic_fsm_stateReg;
  reg        [3:0]    PrivilegedPlugin_logic_fsm_stateNext;
  wire                when_PrivilegedPlugin_l773;
  reg        [2:0]    _zz_PrivilegedPlugin_setup_ramWrite_address;
  reg        [2:0]    _zz_PrivilegedPlugin_setup_ramWrite_address_1;
  reg        [2:0]    _zz_PrivilegedPlugin_setup_ramRead_address;
  reg        [2:0]    _zz_PrivilegedPlugin_setup_ramRead_address_1;
  wire                when_PrivilegedPlugin_l959;
  wire       [1:0]    switch_PrivilegedPlugin_l960;
  wire                when_StateMachine_l253_2;
  `ifndef SYNTHESIS
  reg [31:0] EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string;
  reg [31:0] EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string;
  reg [63:0] ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string;
  reg [39:0] ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [39:0] ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [63:0] ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string;
  reg [31:0] EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string;
  reg [87:0] Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string;
  reg [87:0] Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string;
  reg [31:0] EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string;
  reg [63:0] ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string;
  reg [39:0] ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [39:0] EU0_CsrAccessPlugin_logic_fsm_stateReg_string;
  reg [39:0] EU0_CsrAccessPlugin_logic_fsm_stateNext_string;
  reg [119:0] EnvCallPlugin_logic_flushes_stateReg_string;
  reg [119:0] EnvCallPlugin_logic_flushes_stateNext_string;
  reg [79:0] Lsu2Plugin_logic_special_atomic_stateReg_string;
  reg [79:0] Lsu2Plugin_logic_special_atomic_stateNext_string;
  reg [39:0] MmuPlugin_logic_refill_stateReg_string;
  reg [39:0] MmuPlugin_logic_refill_stateNext_string;
  reg [63:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string;
  reg [63:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string;
  reg [63:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string;
  reg [39:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string;
  reg [39:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string;
  reg [31:0] _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string;
  reg [31:0] _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string;
  reg [31:0] _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string;
  reg [79:0] PrivilegedPlugin_logic_fsm_stateReg_string;
  reg [79:0] PrivilegedPlugin_logic_fsm_stateNext_string;
  `endif

  reg [31:0] FetchCachePlugin_logic_banks_0_mem [0:63];
  (* ram_style = "distributed" *) reg [25:0] FetchCachePlugin_logic_ways_0_mem [0:3];
  (* ram_style = "distributed" *) reg [32:0] BranchContextPlugin_logic_mem_earlyBranch [0:3];
  (* ram_style = "distributed" *) reg [64:0] BranchContextPlugin_logic_mem_finalBranch [0:3];
  (* ram_style = "distributed" *) reg [31:0] DecoderPredictionPlugin_logic_ras_mem_stack [0:15];
  reg [48:0] BtbPlugin_logic_mem [0:7];
  reg [1:0] GSharePlugin_logic_mem_counter [0:127];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_lq_mem_addressPre [0:7];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_lq_mem_addressPost [0:7];
  (* ram_style = "distributed" *) reg [1:0] Lsu2Plugin_logic_lq_mem_size [0:7];
  (* ram_style = "distributed" *) reg [5:0] Lsu2Plugin_logic_lq_mem_physRd [0:7];
  (* ram_style = "distributed" *) reg [3:0] Lsu2Plugin_logic_lq_mem_robId [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_robIdMsb [0:7];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_lq_mem_pc [0:7];
  (* ram_style = "distributed" *) reg [3:0] Lsu2Plugin_logic_lq_mem_sqAlloc [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_io [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_writeRd [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_lr [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_unsigned [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_doSpecial [0:7];
  reg [31:0] Lsu2Plugin_logic_lq_mem_data [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_needTranslation [0:7];
  reg [0:0] Lsu2Plugin_logic_lq_mem_spFpAddress [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_hazardPrediction_valid [0:7];
  (* ram_style = "distributed" *) reg [2:0] Lsu2Plugin_logic_lq_mem_hazardPrediction_delta [0:7];
  (* ram_style = "distributed" *) reg [2:0] Lsu2Plugin_logic_lq_mem_hazardPrediction_score [0:7];
  reg [5:0] Lsu2Plugin_logic_lq_mem_hitPrediction_counter [0:7];
  reg [21:0] Lsu2Plugin_logic_lq_hazardPrediction_mem [0:127];
  reg [5:0] Lsu2Plugin_logic_lq_hitPrediction_mem [0:63];
  (* ram_style = "distributed" *) reg [3:0] Lsu2Plugin_logic_sq_mem_robId [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_robIdMsb [0:7];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_sq_mem_addressPre [0:7];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_sq_mem_addressPost [0:7];
  (* ram_style = "distributed" *) reg [1:0] Lsu2Plugin_logic_sq_mem_size [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_io [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_amo [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_sc [0:7];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_sq_mem_data [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_needTranslation [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_feededOnce [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_doSpecial [0:7];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_doNotBypass [0:7];
  (* ram_style = "distributed" *) reg [3:0] Lsu2Plugin_logic_sq_mem_lqAlloc [0:7];
  (* ram_style = "distributed" *) reg [44:0] FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0 [0:3];
  (* ram_style = "distributed" *) reg [44:0] FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1 [0:3];
  (* ram_style = "distributed" *) reg [44:0] FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2 [0:3];
  (* ram_style = "distributed" *) reg [44:0] FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3 [0:3];
  (* ram_style = "distributed" *) reg [24:0] FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0 [0:3];
  (* ram_style = "distributed" *) reg [24:0] FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1 [0:3];
  (* ram_style = "distributed" *) reg [44:0] Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0 [0:3];
  (* ram_style = "distributed" *) reg [44:0] Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1 [0:3];
  (* ram_style = "distributed" *) reg [44:0] Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2 [0:3];
  (* ram_style = "distributed" *) reg [44:0] Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3 [0:3];
  (* ram_style = "distributed" *) reg [24:0] Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0 [0:3];
  (* ram_style = "distributed" *) reg [24:0] Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1 [0:3];
  (* ram_style = "distributed" *) reg [31:0] CsrRamPlugin_logic_mem [0:7];
  (* ram_style = "distributed" *) reg [26:0] BranchContextPlugin_free_dispatchMem_mem [0:3];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_target [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_1 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_2 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_3 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [31:0] RobPlugin_logic_storage_PC_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_WRITE_RD_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [5:0] RobPlugin_logic_storage_PHYS_RD_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [4:0] RobPlugin_logic_storage_ARCH_RD_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [5:0] RobPlugin_logic_storage_PHYS_RD_FREE_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_BRANCH_SEL_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_BRANCH_TAKEN_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [23:0] RobPlugin_logic_storage_BRANCH_HISTORY_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [3:0] RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_LQ_ALLOC_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_SQ_ALLOC_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [31:0] RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [5:0] RobPlugin_logic_storage_PHYS_RS_0_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_READ_RS_0_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [5:0] RobPlugin_logic_storage_PHYS_RS_1_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_READ_RS_1_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [1:0] RobPlugin_logic_storage_BRANCH_ID_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [3:0] RobPlugin_logic_storage_LSU_ID_banks_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_ROB_MSB_banks_0 [0:15];
  function [31:0] zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue(input dummy);
    begin
      zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue = 32'h00000000;
      zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue[2 : 0] = 3'b101;
    end
  endfunction
  wire [31:0] _zz_259;
  function  zz_DecoderPlugin_logic_slots_0_x0AlwaysZero(input dummy);
    begin
      zz_DecoderPlugin_logic_slots_0_x0AlwaysZero = 1'bx;
      zz_DecoderPlugin_logic_slots_0_x0AlwaysZero = 1'b1;
    end
  endfunction
  wire  _zz_260;

  assign _zz__zz_FetchPlugin_stages_1_MMU_IO = (ioStartAddr + ioSize);
  assign _zz_FetchPlugin_stages_1_FETCH_ID_1 = FetchPlugin_stages_1_isFireing;
  assign _zz_FetchPlugin_stages_1_FETCH_ID = {11'd0, _zz_FetchPlugin_stages_1_FETCH_ID_1};
  assign _zz_FetchCachePlugin_logic_read_onWays_0_hits_bypassHits = (FetchPlugin_stages_1_Fetch_FETCH_PC >>> 4'd8);
  assign _zz_AlignerPlugin_logic_extractors_0_usable = ((_zz_AlignerPlugin_logic_extractors_0_usage ? AlignerPlugin_logic_decoders_0_usable : 1'b0) | (_zz_AlignerPlugin_logic_extractors_0_usage_1 ? AlignerPlugin_logic_decoders_1_usable : 1'b0));
  assign _zz_FrontendPlugin_aligned_PC_0 = (AlignerPlugin_logic_extractors_0_pcWord >>> 2'd2);
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push = (DecoderPredictionPlugin_logic_ras_ptr_push + _zz_DecoderPredictionPlugin_logic_ras_ptr_push_1);
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push_2 = DecoderPredictionPlugin_logic_ras_ptr_pushIt;
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push_1 = {3'd0, _zz_DecoderPredictionPlugin_logic_ras_ptr_push_2};
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push_4 = DecoderPredictionPlugin_logic_ras_ptr_popIt;
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push_3 = {3'd0, _zz_DecoderPredictionPlugin_logic_ras_ptr_push_4};
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop = (DecoderPredictionPlugin_logic_ras_ptr_pop + _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_1);
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_2 = DecoderPredictionPlugin_logic_ras_ptr_pushIt;
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_1 = {3'd0, _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_2};
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_4 = DecoderPredictionPlugin_logic_ras_ptr_popIt;
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_3 = {3'd0, _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_4};
  assign _zz_BtbPlugin_logic_onLearn_port_payload_address = (BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice >>> 2'd2);
  assign _zz_BtbPlugin_logic_readCmd_entryAddress = (FetchPlugin_stages_0_Fetch_FETCH_PC >>> 2'd2);
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_2 = FetchPlugin_stages_0_BRANCH_HISTORY;
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_1 = _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_2[6:0];
  assign _zz_GSharePlugin_logic_onLearn_hash_2 = BranchContextPlugin_free_learn_BRANCH_HISTORY;
  assign _zz_GSharePlugin_logic_onLearn_hash_1 = _zz_GSharePlugin_logic_onLearn_hash_2[6:0];
  assign _zz_CommitPlugin_logic_ptr_allocNext_1 = (FrontendPlugin_allocated_isFireing ? 1'b1 : 1'b0);
  assign _zz_CommitPlugin_logic_ptr_allocNext = {4'd0, _zz_CommitPlugin_logic_ptr_allocNext_1};
  assign _zz_CommitPlugin_logic_reschedule_commit_rowHit = CommitPlugin_logic_ptr_commitRow[3:0];
  assign _zz_CommitPlugin_logic_reschedule_age = CommitPlugin_logic_ptr_free[3:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_0_age = CommitPlugin_logic_ptr_free[3:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_1_age = CommitPlugin_logic_ptr_free[3:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_2_age = CommitPlugin_logic_ptr_free[3:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_3_age = CommitPlugin_logic_ptr_free[3:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_4_age = CommitPlugin_logic_ptr_free[3:0];
  assign _zz_CommitPlugin_logic_reschedule_trap_5 = ((((_zz_CommitPlugin_logic_reschedule_trap ? Lsu2Plugin_setup_sharedTrap_payload_trap : 1'b0) | (_zz_CommitPlugin_logic_reschedule_trap_1 ? 1'b1 : 1'b0)) | ((_zz_CommitPlugin_logic_reschedule_trap_2 ? EU0_BranchPlugin_setup_reschedule_payload_trap : 1'b0) | (_zz_CommitPlugin_logic_reschedule_trap_3 ? 1'b1 : 1'b0))) | (_zz_CommitPlugin_logic_reschedule_trap_4 ? 1'b1 : 1'b0));
  assign _zz_CommitPlugin_logic_reschedule_skipCommit = ((((CommitPlugin_logic_reschedule_portsLogic_hits[0] ? Lsu2Plugin_setup_sharedTrap_payload_skipCommit : 1'b0) | (CommitPlugin_logic_reschedule_portsLogic_hits[1] ? Lsu2Plugin_setup_specialTrap_payload_skipCommit : 1'b0)) | ((CommitPlugin_logic_reschedule_portsLogic_hits[2] ? EU0_BranchPlugin_setup_reschedule_payload_skipCommit : 1'b0) | (CommitPlugin_logic_reschedule_portsLogic_hits[3] ? EnvCallPlugin_setup_reschedule_payload_skipCommit : 1'b0))) | (CommitPlugin_logic_reschedule_portsLogic_hits[4] ? EU0_CsrAccessPlugin_setup_trap_payload_skipCommit : 1'b0));
  assign _zz_CommitPlugin_logic_commit_active_1 = _zz_CommitPlugin_logic_commit_active_2[0 : 0];
  assign _zz_CommitPlugin_logic_commit_active_2 = RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_spinal_port1[0];
  assign _zz_CommitPlugin_logic_commit_head = (CommitPlugin_logic_ptr_commit + 5'h00);
  assign _zz_CommitPlugin_logic_free_robHit = CommitPlugin_logic_ptr_free[3:0];
  assign _zz_commit_pc_0_1 = _zz_commit_pc_0_2[31 : 0];
  assign _zz_commit_pc_0_2 = RobPlugin_logic_storage_PC_banks_0_spinal_port1[31 : 0];
  assign _zz_CommitDebugFilterPlugin_logic_filters_0_value = ($signed(_zz_CommitDebugFilterPlugin_logic_filters_0_value_1) >>> 4);
  assign _zz_CommitDebugFilterPlugin_logic_filters_0_value_1 = _zz_CommitDebugFilterPlugin_logic_filters_0_value_2;
  assign _zz_CommitDebugFilterPlugin_logic_filters_0_value_2 = (_zz_CommitDebugFilterPlugin_logic_filters_0_value_3 - CommitDebugFilterPlugin_logic_filters_0_value);
  assign _zz_CommitDebugFilterPlugin_logic_filters_0_value_3 = {15'd0, CommitDebugFilterPlugin_logic_commits};
  assign _zz_CommitDebugFilterPlugin_logic_filters_1_value = ($signed(_zz_CommitDebugFilterPlugin_logic_filters_1_value_1) >>> 8);
  assign _zz_CommitDebugFilterPlugin_logic_filters_1_value_1 = _zz_CommitDebugFilterPlugin_logic_filters_1_value_2;
  assign _zz_CommitDebugFilterPlugin_logic_filters_1_value_2 = (_zz_CommitDebugFilterPlugin_logic_filters_1_value_3 - CommitDebugFilterPlugin_logic_filters_1_value);
  assign _zz_CommitDebugFilterPlugin_logic_filters_1_value_3 = {15'd0, CommitDebugFilterPlugin_logic_commits};
  assign _zz_CommitDebugFilterPlugin_logic_filters_2_value = ($signed(_zz_CommitDebugFilterPlugin_logic_filters_2_value_1) >>> 12);
  assign _zz_CommitDebugFilterPlugin_logic_filters_2_value_1 = _zz_CommitDebugFilterPlugin_logic_filters_2_value_2;
  assign _zz_CommitDebugFilterPlugin_logic_filters_2_value_2 = (_zz_CommitDebugFilterPlugin_logic_filters_2_value_3 - CommitDebugFilterPlugin_logic_filters_2_value);
  assign _zz_CommitDebugFilterPlugin_logic_filters_2_value_3 = {15'd0, CommitDebugFilterPlugin_logic_commits};
  assign _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_1 = _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_2[31 : 0];
  assign _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_2 = RobPlugin_logic_storage_PC_banks_0_spinal_port2[31 : 0];
  assign _zz__zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1) + $signed(ALU0_SrcPlugin_logic_addsub_rs2Patched));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1 = _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2 = {31'd0, _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3};
  assign _zz_ALU0_IntAluPlugin_logic_process_result_1 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
  assign _zz_ALU0_IntAluPlugin_logic_process_result = {31'd0, _zz_ALU0_IntAluPlugin_logic_process_result_1};
  assign _zz_ALU0_ShiftPlugin_logic_process_amplitude = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[4 : 0];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed = {ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[0],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[1],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[2],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[3],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[4],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[5],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[6],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[7],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[8],{_zz_ALU0_ShiftPlugin_logic_process_reversed_1,{_zz_ALU0_ShiftPlugin_logic_process_reversed_2,_zz_ALU0_ShiftPlugin_logic_process_reversed_3}}}}}}}}}}};
  assign _zz_ALU0_ShiftPlugin_logic_process_shifted = ($signed(_zz_ALU0_ShiftPlugin_logic_process_shifted_1) >>> ALU0_ShiftPlugin_logic_process_amplitude);
  assign _zz_ALU0_ShiftPlugin_logic_process_shifted_1 = {(ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED && ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]),ALU0_ShiftPlugin_logic_process_reversed};
  assign _zz_ALU0_ShiftPlugin_logic_process_patched = {ALU0_ShiftPlugin_logic_process_shifted[0],{ALU0_ShiftPlugin_logic_process_shifted[1],{ALU0_ShiftPlugin_logic_process_shifted[2],{ALU0_ShiftPlugin_logic_process_shifted[3],{ALU0_ShiftPlugin_logic_process_shifted[4],{ALU0_ShiftPlugin_logic_process_shifted[5],{ALU0_ShiftPlugin_logic_process_shifted[6],{ALU0_ShiftPlugin_logic_process_shifted[7],{ALU0_ShiftPlugin_logic_process_shifted[8],{_zz_ALU0_ShiftPlugin_logic_process_patched_1,{_zz_ALU0_ShiftPlugin_logic_process_patched_2,_zz_ALU0_ShiftPlugin_logic_process_patched_3}}}}}}}}}}};
  assign _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 25],EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[11 : 7]};
  assign _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2_1 = EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1) + $signed(EU0_SrcPlugin_logic_addsub_rs2Patched));
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3 = EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2 = {31'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED_1 = EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED = {31'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED_1 = EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED = {31'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[0] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2 = {{31{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[1] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4 = {{30{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[2] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6 = {{29{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[3] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8 = {{28{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[4] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10 = {{27{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[5] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12 = {{26{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[6] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14 = {{25{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[7] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16 = {{24{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[8] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18 = {{23{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[9] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20 = {{22{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[10] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22 = {{21{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[11] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24 = {{20{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[12] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26 = {{19{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[13] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28 = {{18{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[14] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30 = {{17{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[15] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32 = {{16{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[16] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34 = {{15{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[17] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36 = {{14{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[18] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38 = {{13{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[19] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40 = {{12{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[20] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42 = {{11{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[21] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44 = {{10{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[22] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46 = {{9{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[23] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48 = {{8{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[24] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50 = {{7{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[25] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52 = {{6{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[26] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54 = {{5{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[27] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56 = {{4{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[28] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58 = {{3{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[29] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60 = {{2{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[30] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62 = {{1{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62_1[0]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_63 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[31] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 32] : 1'b0);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_1 = ($signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_2) * $signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_3));
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_1[31:0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_2 = {1'b0,EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0]};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64_3 = EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[32 : 32];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_5 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_6);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_9);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_8 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_9 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_12);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_9 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_10 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_11 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_12 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_13 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_14);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_14 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_19);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_16 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_17 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_19 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_20 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_21);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_20 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_21 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_12);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_9 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_10 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_11 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_12 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_13 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_14);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_14 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_19);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_16 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_17 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_19 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_20 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_21);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_20 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_21 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_12);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_9 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_10 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_11 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_12 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_13 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_14);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_14 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_19);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_16 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_17 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_19 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_20 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_21);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_20 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_21 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_12);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_9 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_10 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_11 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_12 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_13 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_14);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_14 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_19);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_16 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_17 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_19 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_20 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_21);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_20 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_21 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_12);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_9 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_10 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_11 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_12 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_13 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_14);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_14 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_19);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_16 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_17 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_19 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_20 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_21);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_20 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_21 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_12);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_9 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_10 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_11 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_12 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_13 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_14);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_14 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_19);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_16 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_17 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_19 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_20 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_21);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_20 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_21 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_12);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_9 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_10 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_11 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_12 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_13 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_14);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_14 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_19);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_16 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_17 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_19 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_20 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_21);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_20 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_21 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_12);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_9 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_10 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_11 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_12 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_13 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_14);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_14 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_19);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_16 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_17 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_19 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_20 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_21);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_20 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_6};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_21 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_7};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_11);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_9 + _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_10);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_9 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_10 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_11 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_12 + _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_13);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_12 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_13 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_14 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_15 + _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_18);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_15 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_16 + _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_17);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_16 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_4};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_17 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_5};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_18 = {3'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_6};
  assign _zz_EU0_DivPlugin_logic_rsp_selected = {2'd0, EU0_DivPlugin_logic_div_io_rsp_payload_remain};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_1 = _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_2;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_2 = ((EU0_ExecutionUnitBase_pipeline_execute_1_DIV_REVERT_RESULT ? (~ _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT) : _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT) + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_3);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_4 = EU0_ExecutionUnitBase_pipeline_execute_1_DIV_REVERT_RESULT;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_3 = {34'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_4};
  assign _zz_EU0_BranchPlugin_logic_process_target_b = {{{{EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31],EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[19 : 12]},EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[20]},EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[30 : 21]},1'b0};
  assign _zz_EU0_BranchPlugin_logic_process_target_b_1 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_EU0_BranchPlugin_logic_process_target_b_2 = {{{{EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31],EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[7]},EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[30 : 25]},EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[11 : 8]},1'b0};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE = ($signed(EU0_BranchPlugin_logic_process_target_a) + $signed(EU0_BranchPlugin_logic_process_target_b));
  assign _zz_EU0_BranchPlugin_logic_process_slices_1 = 1'b0;
  assign _zz_EU0_BranchPlugin_logic_process_slices = {1'd0, _zz_EU0_BranchPlugin_logic_process_slices_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1 = ({2'd0,EU0_BranchPlugin_logic_process_slices} <<< 2'd2);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE = {28'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1};
  assign _zz_LsuPlugin_peripheralBus_toAxiLite4_addr = ({2'd0,LsuPlugin_peripheralBus_toAxiLite4_a_payload_address[31 : 2]} <<< 2'd2);
  assign _zz_BranchContextPlugin_logic_onCommit_commitedNext = {2'd0, _zz_BranchContextPlugin_logic_onCommit_commitedNext_1};
  assign _zz_HistoryPlugin_logic_onCommit_valueNext_1 = {HistoryPlugin_logic_onCommit_valueNext,HistoryPlugin_logic_onCommit_isTaken_0};
  assign _zz_HistoryPlugin_logic_update_pushes_0_stateNext_1 = {HistoryPlugin_logic_update_pushes_0_stateNext,BtbPlugin_setup_historyPush_taken[0]};
  assign _zz_HistoryPlugin_logic_update_pushes_2_stateNext_1 = {HistoryPlugin_logic_update_pushes_2_stateNext,DecoderPredictionPlugin_setup_historyPush_taken[0]};
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_1 = _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_2[23 : 0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_2 = RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_spinal_port1[23 : 0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_1 = _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_2[0 : 0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_2 = RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_spinal_port2[0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_1 = _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_2[0 : 0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_2 = RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_spinal_port2[0];
  assign _zz_DecoderPredictionPlugin_logic_ras_healPush_1 = _zz_DecoderPredictionPlugin_logic_ras_healPush_2[3 : 0];
  assign _zz_DecoderPredictionPlugin_logic_ras_healPush_2 = RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_spinal_port1[3 : 0];
  assign _zz_Lsu2Plugin_logic_lq_tracker_freeNext = (Lsu2Plugin_logic_lq_tracker_free + _zz_Lsu2Plugin_logic_lq_tracker_freeNext_1);
  assign _zz_Lsu2Plugin_logic_lq_tracker_freeNext_1 = {3'd0, Lsu2Plugin_logic_lq_tracker_add};
  assign _zz_Lsu2Plugin_logic_lq_tracker_freeNext_2 = {3'd0, Lsu2Plugin_logic_lq_tracker_sub};
  assign _zz_when_Lsu2Plugin_l454 = Lsu2Plugin_logic_lq_onCommit_free[2:0];
  assign _zz_when_Lsu2Plugin_l454_1 = Lsu2Plugin_logic_lq_onCommit_free[2:0];
  assign _zz_when_Lsu2Plugin_l454_2 = Lsu2Plugin_logic_lq_onCommit_free[2:0];
  assign _zz_when_Lsu2Plugin_l454_3 = Lsu2Plugin_logic_lq_onCommit_free[2:0];
  assign _zz_when_Lsu2Plugin_l454_4 = Lsu2Plugin_logic_lq_onCommit_free[2:0];
  assign _zz_when_Lsu2Plugin_l454_5 = Lsu2Plugin_logic_lq_onCommit_free[2:0];
  assign _zz_when_Lsu2Plugin_l454_6 = Lsu2Plugin_logic_lq_onCommit_free[2:0];
  assign _zz_when_Lsu2Plugin_l454_7 = Lsu2Plugin_logic_lq_onCommit_free[2:0];
  assign _zz_Lsu2Plugin_logic_lq_onCommit_priority_1 = (Lsu2Plugin_logic_lq_onCommit_priority <<< 1);
  assign _zz_Lsu2Plugin_logic_lq_onCommit_free_1_1 = Lsu2Plugin_logic_lq_onCommit_lqCommits_0;
  assign _zz_Lsu2Plugin_logic_lq_onCommit_free_1 = {3'd0, _zz_Lsu2Plugin_logic_lq_onCommit_free_1_1};
  assign _zz_Lsu2Plugin_logic_lq_ptr_free = {3'd0, Lsu2Plugin_logic_lq_onCommit_lqCommitCount};
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext = (_zz_Lsu2Plugin_logic_sq_tracker_freeNext_1 - _zz_Lsu2Plugin_logic_sq_tracker_freeNext_3);
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext_1 = (_zz_Lsu2Plugin_logic_sq_tracker_freeNext_2 - Lsu2Plugin_logic_sq_ptr_alloc);
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext_2 = (4'b1000 + Lsu2Plugin_logic_sq_ptr_free);
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext_3 = {3'd0, Lsu2Plugin_logic_sq_tracker_sub};
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext_4 = {3'd0, Lsu2Plugin_logic_sq_tracker_add};
  assign _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1_1 = when_Lsu2Plugin_l591;
  assign _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1 = {3'd0, _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1_1};
  assign _zz_Lsu2Plugin_logic_lq_mem_addressPre_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_physRd_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_robId_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_pc_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_writeRd_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_lr_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_size_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_unsigned_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_needTranslation_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPre_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_robId_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_amo_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_sc_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_size_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_needTranslation_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_data_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh = ({1'd0,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pHigh} <<< 1'd1);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh = ({1'd0,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pHigh} <<< 1'd1);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s1_cmp = (Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ROB_FULL - Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ROB_FULL);
  assign _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu = ({AguPlugin_setup_port_payload_robIdMsb,AguPlugin_setup_port_payload_robId} - Lsu2Plugin_logic_sharedPip_stages_0_LQ_ROB_FULL);
  assign _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu_1 = ({AguPlugin_setup_port_payload_robIdMsb,AguPlugin_setup_port_payload_robId} - Lsu2Plugin_logic_sharedPip_stages_0_SQ_ROB_FULL);
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID = ((Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ || (! Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask)) ? Lsu2Plugin_logic_sharedPip_stages_0_LQ_ROB_FULL : Lsu2Plugin_logic_sharedPip_stages_0_SQ_ROB_FULL);
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_1 = {AguPlugin_setup_port_payload_robIdMsb,AguPlugin_setup_port_payload_robId};
  assign _zz_Lsu2Plugin_logic_lq_mem_sqAlloc_port_1 = _zz_Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC[2:0];
  assign _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT = (Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC - _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1);
  assign _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1 = {1'd0, Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1 = (_zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT - Lsu2Plugin_logic_sq_ptr_free);
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh = {1'd0, Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pLow};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh = ({1'd0,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pHigh} <<< 1'd1);
  assign _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta = (_zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_1 - 4'b0001);
  assign _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_1 = (Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port4 - _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_2);
  assign _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_2 = {1'd0, Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID};
  assign _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_1 = {Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION_COUNTER[5],Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION_COUNTER};
  assign _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_2 = {_zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[5],_zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next};
  assign _zz_when_SInt_l132 = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[6 : 5];
  assign _zz_when_SInt_l138 = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[5 : 5];
  assign _zz_Lsu2Plugin_logic_sq_ptr_writeBack_1 = Lsu2Plugin_logic_writeback_feed_fire;
  assign _zz_Lsu2Plugin_logic_sq_ptr_writeBack = {3'd0, _zz_Lsu2Plugin_logic_sq_ptr_writeBack_1};
  assign _zz_Lsu2Plugin_setup_specialTrap_payload_cause = (Lsu2Plugin_logic_special_isStore ? 3'b111 : 3'b101);
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_2 = ($signed(_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_3) + $signed(_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_6));
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_3 = ($signed(_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_4) + $signed(_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_5));
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_4 = _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1;
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_5 = (Lsu2Plugin_logic_special_atomic_alu_compare ? (~ _zz_Lsu2Plugin_logic_special_atomic_alu_addSub) : _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_7 = (Lsu2Plugin_logic_special_atomic_alu_compare ? 2'b01 : 2'b00);
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_6 = {{30{_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_7[1]}}, _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_7};
  assign _zz_EU0_BranchPlugin_setup_intFormatPort_payload = EU0_ExecutionUnitBase_pipeline_execute_2_PC_FALSE;
  assign _zz_EU0_BranchPlugin_setup_reschedule_payload_reason = ((EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL == BranchPlugin_BranchCtrlEnum_B) ? 5'h10 : 5'h11);
  assign _zz_EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1 = 2'b00;
  assign _zz_EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice = {30'd0, _zz_EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement;
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext = {1'd0, _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement;
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext = {1'd0, _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_6 = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowExecute : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowExecute : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowExecute : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowExecute : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowExecute : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowExecute : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowRead : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowRead : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowRead : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowRead : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowRead : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowRead : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowWrite : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowWrite : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowWrite : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowWrite : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowWrite : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowWrite : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowUser : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowUser : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowUser : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowUser : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowUser : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowUser : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_pageFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_pageFault : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_pageFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_pageFault : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_pageFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_pageFault : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_accessFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_accessFault : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_accessFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_accessFault : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_accessFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_accessFault : 1'b0)));
  assign _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input - 3'b001);
  assign _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input - 2'b01);
  assign _zz_EU0_CsrAccessPlugin_setup_onDecodeAddress = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
  assign _zz_EU0_CsrAccessPlugin_setup_onReadAddress = EU0_CsrAccessPlugin_logic_fsm_regs_microOp;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1 = EU0_CsrAccessPlugin_logic_fsm_regs_microOp[19 : 15];
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = {27'd0, _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1};
  assign _zz_EU0_CsrAccessPlugin_setup_onWriteAddress = EU0_CsrAccessPlugin_logic_fsm_regs_microOp;
  assign _zz_csrAccess_payload_address = EU0_ExecutionUnitBase_pipeline_execute_2_Frontend_MICRO_OP;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_6 = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowExecute : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowExecute : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowExecute : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowExecute : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowExecute : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowExecute : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowRead : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowRead : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowRead : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowRead : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowRead : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowRead : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowWrite : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowWrite : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowWrite : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowWrite : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowWrite : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowWrite : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowUser : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowUser : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowUser : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowUser : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowUser : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowUser : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineException = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_pageFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_pageFault : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_pageFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_pageFault : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_pageFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_pageFault : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_accessFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_accessFault : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_accessFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_accessFault : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_accessFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_accessFault : 1'b0)));
  assign _zz_MmuPlugin_logic_refill_portsRequests_ohFirst_masked = (MmuPlugin_logic_refill_portsRequests_ohFirst_input - 2'b01);
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask_1 = (4'b0001 <<< FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value);
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask_1 = (4'b0001 <<< Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value);
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask = (2'b01 <<< FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value);
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask = (2'b01 <<< Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value);
  assign _zz_FrontendPlugin_decoded_READ_RS_0_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000044) == 32'h00000000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000018) == 32'h00000000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00006004) == 32'h00002000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00005004) == 32'h00001000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00002050) == 32'h00002000)}}}});
  assign _zz_FrontendPlugin_decoded_READ_RS_1_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000034) == 32'h00000020),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000064) == 32'h00000020),{_zz_FrontendPlugin_decoded_SQ_ALLOC_0_1,_zz_FrontendPlugin_decoded_SQ_ALLOC_0}}});
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_1 = (|{_zz_FrontendPlugin_decoded_WRITE_RD_0,{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00001010) == 32'h00001010),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00002010) == 32'h00002010),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_WRITE_RD_0_2) == 32'h00002008),{(_zz_FrontendPlugin_decoded_WRITE_RD_0_3 == _zz_FrontendPlugin_decoded_WRITE_RD_0_4),{_zz_FrontendPlugin_decoded_WRITE_RD_0_5,_zz_FrontendPlugin_decoded_WRITE_RD_0_6}}}}}});
  assign _zz_FrontendPlugin_decoded_ALU0_SEL_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000030) == 32'h00000010),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000004c) == 32'h00000004),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h02000050) == 32'h00000010)}});
  assign _zz_FrontendPlugin_decoded_EU0_SEL_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000040) == 32'h00000040),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000010) == 32'h00000000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h02000024) == 32'h02000020)}});
  assign _zz_FrontendPlugin_decoded_LQ_ALLOC_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000038) == 32'h00000000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h18002048) == 32'h10002008)});
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_0_2 = (|{_zz_FrontendPlugin_decoded_SQ_ALLOC_0_1,{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000078) == 32'h00000020),_zz_FrontendPlugin_decoded_SQ_ALLOC_0}});
  assign _zz_DecoderPlugin_logic_exception_compressedFault = (DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_compressedFaultReg_0 : 1'b0);
  assign _zz_DecoderPlugin_logic_exception_fetchFault = (DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_fetchFaultReg_0 : 1'b0);
  assign _zz_DecoderPlugin_logic_exception_fetchFaultPage = (DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_fetchFaultPageReg_0 : 1'b0);
  assign _zz_DecoderPlugin_logic_exception_debugEnter = (DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_debugEnterReg_0 : 1'b0);
  assign _zz_DecoderPlugin_setup_exceptionPort_payload_tval = (DecoderPlugin_logic_exception_pc + _zz_DecoderPlugin_setup_exceptionPort_payload_tval_1);
  assign _zz_DecoderPlugin_setup_exceptionPort_payload_tval_2 = 2'b00;
  assign _zz_DecoderPlugin_setup_exceptionPort_payload_tval_1 = {30'd0, _zz_DecoderPlugin_setup_exceptionPort_payload_tval_2};
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_1[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_1 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_3,{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_2,{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0,((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h10002048) == 32'h10002008)}}}});
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_1[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_1 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_3,{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_1,{((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h08002048) == 32'h08002008),((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h10002048) == 32'h00002008)}}});
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_4 = _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_5[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_5 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_3,{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_2,{_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_1,{((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h00002048) == 32'h00002008),_zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0}}}});
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0_1[0];
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0_1 = 1'b0;
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0_1[0];
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0_1 = 1'b0;
  assign _zz_FrontendPlugin_decoded_OP_ID_1 = FrontendPlugin_decoded_isFireing;
  assign _zz_FrontendPlugin_decoded_OP_ID = {11'd0, _zz_FrontendPlugin_decoded_OP_ID_1};
  assign _zz_FrontendPlugin_decoded_IS_JAL_0 = (|_zz_FrontendPlugin_decoded_WRITE_RD_0);
  assign _zz_FrontendPlugin_decoded_IS_JALR_0 = (|((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000001c) == 32'h00000004));
  assign _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_0 = (|((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000054) == 32'h00000040));
  assign _zz_FrontendPlugin_decoded_IS_ANY_0 = (|((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000050) == 32'h00000040));
  assign _zz__zz_FrontendPlugin_decoded_OFFSET_0 = {{{{FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[31],FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[7]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[30 : 25]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[11 : 8]},1'b0};
  assign _zz__zz_FrontendPlugin_decoded_OFFSET_0_1 = {{{{FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[31],FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[19 : 12]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[20]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[30 : 21]},1'b0};
  assign _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices_1 = 1'b0;
  assign _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices = {1'd0, _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices_1};
  assign _zz_FrontendPlugin_decoded_PC_INC_0 = (FrontendPlugin_decoded_PC_0 + _zz_FrontendPlugin_decoded_PC_INC_0_1);
  assign _zz_FrontendPlugin_decoded_PC_INC_0_2 = ({2'd0,DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices} <<< 2'd2);
  assign _zz_FrontendPlugin_decoded_PC_INC_0_1 = {28'd0, _zz_FrontendPlugin_decoded_PC_INC_0_2};
  assign _zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0 = FrontendPlugin_decoded_PC_0;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2 = RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_spinal_port1[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2[5 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2 = RobPlugin_logic_storage_PHYS_RS_0_banks_0_spinal_port1[5 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2[0 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2 = RobPlugin_logic_storage_READ_RS_0_banks_0_spinal_port1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2[5 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2 = RobPlugin_logic_storage_PHYS_RS_1_banks_0_spinal_port1[5 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2[0 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2 = RobPlugin_logic_storage_READ_RS_1_banks_0_spinal_port1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2[0 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2 = RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port3[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_2[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_2 = RobPlugin_logic_storage_PC_banks_0_spinal_port3[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2 = (|{((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002000) == 32'h00002000),{_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL,((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001000) == 32'h00000000)}});
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000000) == 32'h00000000));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00003004) == 32'h00001000));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004000) == 32'h00000000));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h40000000) == 32'h40000000));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1 = (|{((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002004) == 32'h00002000),((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h40000024) == 32'h40000020)});
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000024) == 32'h00000024));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_2[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_2 = (|_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2[31 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2 = RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_spinal_port2[31 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2 = RobPlugin_logic_storage_READ_RS_0_banks_0_spinal_port2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2 = RobPlugin_logic_storage_READ_RS_1_banks_0_spinal_port2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2 = RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port4[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_2[31 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_2 = RobPlugin_logic_storage_PC_banks_0_spinal_port4[31 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2[1 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2 = RobPlugin_logic_storage_BRANCH_ID_banks_0_spinal_port1[1 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_2[3 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_2 = RobPlugin_logic_storage_LSU_ID_banks_0_spinal_port1[3 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_2[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_2 = RobPlugin_logic_storage_ROB_MSB_banks_0_spinal_port1[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004050) == 32'h00000010));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2_1 = (|{_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT,{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000010) == 32'h00000010),((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002008) == 32'h00000008)}});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH_1 = (|{_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR,_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED_1 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001000) == 32'h00000000),_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_2 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00005000) == 32'h00004000),_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004060) == 32'h00004020));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM_1 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000050) == 32'h00000040));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL_1 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002050) == 32'h00002000),((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000058) == 32'h00000000)});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h10000008) == 32'h00000008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h10000008) == 32'h10000008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_2 = (|{_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD,((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h18000008) == 32'h10000008)});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT_1 = 1'b0;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000020) == 32'h00000020));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h12103010) == 32'h00000010));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h12103010) == 32'h00100010));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h12403010) == 32'h10000010));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h12203010) == 32'h10000010));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00003048) == 32'h00000008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00005048) == 32'h00001008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h12003010) == 32'h12000010));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004048) == 32'h00004008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL_1 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001050) == 32'h00001050),((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002050) == 32'h00002050)});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004000) == 32'h00004000));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_1 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_2 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_2 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_2 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED);
  assign _zz_BranchContextPlugin_free_learn_GSHARE_COUNTER_0 = BranchContextPlugin_free_learn_raw[25 : 24];
  assign _zz_DispatchPlugin_logic_ptr_next = (CommitPlugin_logic_commit_reschedulePort_payload_robIdNext - 4'b1000);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_0 = (8'h01 <<< _zz_DispatchPlugin_logic_push_slots_0_events_0_1);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_0_2 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0 - DispatchPlugin_logic_ptr_next);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_0_1 = _zz_DispatchPlugin_logic_push_slots_0_events_0_2[2:0];
  assign _zz_DispatchPlugin_logic_push_slots_0_events_1 = (8'h01 <<< _zz_DispatchPlugin_logic_push_slots_0_events_1_1);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_1_2 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0 - DispatchPlugin_logic_ptr_next);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_1_1 = _zz_DispatchPlugin_logic_push_slots_0_events_1_2[2:0];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID = {1'd0, DispatchPlugin_logic_pop_0_stagesList_1_UINT};
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID = {1'd0, DispatchPlugin_logic_pop_1_stagesList_1_UINT};
  assign _zz_DispatchPlugin_logic_wake_dynamic_offseted_0_payload = (Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_payload_robId - DispatchPlugin_logic_ptr_current);
  assign _zz_DispatchPlugin_logic_wake_dynamic_offseted_1_payload = (Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_payload_robId - DispatchPlugin_logic_ptr_current);
  assign _zz_DispatchPlugin_logic_wake_dynamic_offseted_2_payload = (Lsu2Plugin_logic_special_wakeRob_payload_robId - DispatchPlugin_logic_ptr_current);
  assign _zz_DispatchPlugin_logic_wake_dynamic_offseted_3_payload = (EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_payload_robId - DispatchPlugin_logic_ptr_current);
  assign _zz_DispatchPlugin_logic_wake_dynamic_masks_0 = (8'h01 <<< DispatchPlugin_logic_wake_dynamic_offseted_0_payload);
  assign _zz_DispatchPlugin_logic_wake_dynamic_masks_1 = (8'h01 <<< DispatchPlugin_logic_wake_dynamic_offseted_1_payload);
  assign _zz_DispatchPlugin_logic_wake_dynamic_masks_2 = (8'h01 <<< DispatchPlugin_logic_wake_dynamic_offseted_2_payload);
  assign _zz_DispatchPlugin_logic_wake_dynamic_masks_3 = (8'h01 <<< DispatchPlugin_logic_wake_dynamic_offseted_3_payload);
  assign _zz_integer_RfAllocationPlugin_logic_push_mask_0_1 = _zz_integer_RfAllocationPlugin_logic_push_mask_0_2[0 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_mask_0_2 = RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_spinal_port2[0];
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1 = _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_2[0 : 0];
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_2 = RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port1[0];
  assign _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1 = _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_2[0 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_2 = RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port2[0];
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_1 = _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2[5 : 0];
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2 = RobPlugin_logic_storage_PHYS_RD_banks_0_spinal_port1[5 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_1 = _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2[5 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2 = RobPlugin_logic_storage_PHYS_RD_banks_0_spinal_port2[5 : 0];
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_1 = _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2[4 : 0];
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2 = RobPlugin_logic_storage_ARCH_RD_banks_0_spinal_port1[4 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_1 = _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2[5 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2 = RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_spinal_port1[5 : 0];
  assign _zz_BranchContextPlugin_logic_onCommit_isBranch_0_1 = _zz_BranchContextPlugin_logic_onCommit_isBranch_0_2[0 : 0];
  assign _zz_BranchContextPlugin_logic_onCommit_isBranch_0_2 = RobPlugin_logic_storage_BRANCH_SEL_banks_0_spinal_port1[0];
  assign _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1 = _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_2[0 : 0];
  assign _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_2 = RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_spinal_port1[0];
  assign _zz_HistoryPlugin_logic_onCommit_isTaken_0_1 = _zz_HistoryPlugin_logic_onCommit_isTaken_0_2[0 : 0];
  assign _zz_HistoryPlugin_logic_onCommit_isTaken_0_2 = RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_spinal_port1[0];
  assign _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_1 = _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2[0 : 0];
  assign _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2 = RobPlugin_logic_storage_LQ_ALLOC_banks_0_spinal_port1[0];
  assign _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_1 = _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2[0 : 0];
  assign _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2 = RobPlugin_logic_storage_SQ_ALLOC_banks_0_spinal_port1[0];
  assign _zz_PcPlugin_logic_init_counter_1 = (! PcPlugin_logic_init_booted);
  assign _zz_PcPlugin_logic_init_counter = {6'd0, _zz_PcPlugin_logic_init_counter_1};
  assign _zz_PcPlugin_logic_fetchPc_pc_1 = ({2'd0,PcPlugin_logic_fetchPc_inc} <<< 2'd2);
  assign _zz_PcPlugin_logic_fetchPc_pc = {29'd0, _zz_PcPlugin_logic_fetchPc_pc_1};
  assign _zz_PrivilegedPlugin_setup_ramWrite_data = PrivilegedPlugin_logic_reschedule_payload_epc;
  assign _zz_PrivilegedPlugin_setup_ramWrite_data_1 = PrivilegedPlugin_logic_reschedule_payload_tval;
  assign _zz_PrivilegedPlugin_logic_readed = (PrivilegedPlugin_logic_reschedule_payload_epc + _zz_PrivilegedPlugin_logic_readed_1);
  assign _zz_PrivilegedPlugin_logic_readed_2 = ((PrivilegedPlugin_logic_reschedule_payload_cause != 4'b1010) ? _zz_PrivilegedPlugin_logic_readed_3 : 4'b0000);
  assign _zz_PrivilegedPlugin_logic_readed_1 = {28'd0, _zz_PrivilegedPlugin_logic_readed_2};
  assign _zz_PrivilegedPlugin_logic_readed_3 = ({2'd0,_zz_PrivilegedPlugin_logic_readed_4} <<< 2'd2);
  assign _zz_PrivilegedPlugin_logic_readed_4 = (_zz_PrivilegedPlugin_logic_readed_5 + {1'b0,1'b1});
  assign _zz_PrivilegedPlugin_logic_readed_6 = 1'b0;
  assign _zz_PrivilegedPlugin_logic_readed_5 = {1'd0, _zz_PrivilegedPlugin_logic_readed_6};
  assign _zz_FetchCachePlugin_logic_ways_0_mem_port = {FetchCachePlugin_logic_waysWrite_tag_address,{FetchCachePlugin_logic_waysWrite_tag_error,FetchCachePlugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchCachePlugin_logic_ways_0_mem_port_1 = FetchCachePlugin_logic_waysWrite_mask[0];
  assign _zz_BranchContextPlugin_logic_mem_earlyBranch_port = {FrontendPlugin_allocated_BRANCH_EARLY_0_pc,FrontendPlugin_allocated_BRANCH_EARLY_0_taken};
  assign _zz_BranchContextPlugin_logic_mem_finalBranch_port = {EU0_BranchPlugin_logic_branch_finalBranch_payload_data_taken,{EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget,EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice}};
  assign _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port = DecoderPredictionPlugin_logic_ras_write_payload_data;
  assign _zz_BtbPlugin_logic_mem_port = {BtbPlugin_logic_onLearn_port_payload_data_isBranch,{BtbPlugin_logic_onLearn_port_payload_data_pcTarget,BtbPlugin_logic_onLearn_port_payload_data_hash}};
  assign _zz_GSharePlugin_logic_mem_counter_port = GSharePlugin_logic_mem_write_payload_data_0;
  assign _zz_Lsu2Plugin_logic_lq_mem_addressPre_port_1 = AguPlugin_setup_port_payload_address;
  assign _zz_Lsu2Plugin_logic_lq_mem_addressPost_port = Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
  assign _zz_Lsu2Plugin_logic_lq_mem_size_port_1 = AguPlugin_setup_port_payload_size;
  assign _zz_Lsu2Plugin_logic_lq_mem_physRd_port_1 = AguPlugin_setup_port_payload_physicalRd;
  assign _zz_Lsu2Plugin_logic_lq_mem_robId_port_1 = AguPlugin_setup_port_payload_robId;
  assign _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port_1 = AguPlugin_setup_port_payload_robIdMsb;
  assign _zz_Lsu2Plugin_logic_lq_mem_pc_port_1 = AguPlugin_setup_port_payload_pc;
  assign _zz_Lsu2Plugin_logic_lq_mem_sqAlloc_port = Lsu2Plugin_logic_allocation_stores_alloc;
  assign _zz_Lsu2Plugin_logic_lq_mem_io_port = Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO;
  assign _zz_Lsu2Plugin_logic_lq_mem_writeRd_port_1 = AguPlugin_setup_port_payload_writeRd;
  assign _zz_Lsu2Plugin_logic_lq_mem_lr_port_1 = AguPlugin_setup_port_payload_lr;
  assign _zz_Lsu2Plugin_logic_lq_mem_unsigned_port_1 = AguPlugin_setup_port_payload_unsigned;
  assign _zz_Lsu2Plugin_logic_lq_mem_doSpecial_port = 1'b0;
  assign _zz_Lsu2Plugin_logic_lq_mem_doSpecial_port_1 = 1'b1;
  assign _zz_Lsu2Plugin_logic_lq_mem_needTranslation_port_1 = 1'b1;
  assign _zz_Lsu2Plugin_logic_lq_mem_needTranslation_port_2 = Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO;
  assign _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port = (|{(FrontendPlugin_dispatch_ARCH_RS_0_0 == 5'h08),{(FrontendPlugin_dispatch_ARCH_RS_0_0 == 5'h03),(FrontendPlugin_dispatch_ARCH_RS_0_0 == 5'h02)}});
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port_1 = Lsu2Plugin_logic_aguPush_0_hazardPrediction_hit;
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port_1 = Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_delta;
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port_1 = Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
  assign _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port_1 = Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
  assign _zz_Lsu2Plugin_logic_lq_hazardPrediction_mem_port = {Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_delta,{Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_tag,Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_score}};
  assign _zz_Lsu2Plugin_logic_lq_hitPrediction_mem_port = Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_data_counter;
  assign _zz_Lsu2Plugin_logic_sq_mem_robId_port_1 = AguPlugin_setup_port_payload_robId;
  assign _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port_1 = AguPlugin_setup_port_payload_robIdMsb;
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPre_port_1 = AguPlugin_setup_port_payload_address;
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPost_port = Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
  assign _zz_Lsu2Plugin_logic_sq_mem_size_port_1 = AguPlugin_setup_port_payload_size;
  assign _zz_Lsu2Plugin_logic_sq_mem_io_port = Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO;
  assign _zz_Lsu2Plugin_logic_sq_mem_amo_port_1 = AguPlugin_setup_port_payload_amo;
  assign _zz_Lsu2Plugin_logic_sq_mem_sc_port_1 = AguPlugin_setup_port_payload_sc;
  assign _zz_Lsu2Plugin_logic_sq_mem_needTranslation_port_1 = 1'b1;
  assign _zz_Lsu2Plugin_logic_sq_mem_needTranslation_port_2 = Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO;
  assign _zz_Lsu2Plugin_logic_sq_mem_feededOnce_port = 1'b0;
  assign _zz_Lsu2Plugin_logic_sq_mem_feededOnce_port_1 = 1'b1;
  assign _zz_Lsu2Plugin_logic_sq_mem_doSpecial_port = 1'b0;
  assign _zz_Lsu2Plugin_logic_sq_mem_doSpecial_port_1 = 1'b1;
  assign _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port_1 = (AguPlugin_setup_port_payload_amo || AguPlugin_setup_port_payload_sc);
  assign _zz_Lsu2Plugin_logic_sq_mem_lqAlloc_port = Lsu2Plugin_logic_allocation_loads_alloc_1;
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port = {FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask[0];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port = {FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask[1];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port = {FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask[2];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port = {FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask[3];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port = {FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask[0];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port = {FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask[1];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port = {Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask[0];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port = {Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask[1];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port = {Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask[2];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port = {Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask[3];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port = {Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask[0];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port = {Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask[1];
  assign _zz_RobPlugin_logic_completionMem_hits_0_port = (! RobPlugin_logic_completionMem_hits_0_spinal_port1[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_1_port = (! RobPlugin_logic_completionMem_hits_1_spinal_port1[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_2_port = (! RobPlugin_logic_completionMem_hits_2_spinal_port1[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_3_port = (! RobPlugin_logic_completionMem_hits_3_spinal_port1[0]);
  assign _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port = FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0;
  assign _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PC_banks_0_port = FrontendPlugin_allocated_PC_0;
  assign _zz_RobPlugin_logic_storage_PC_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port = FrontendPlugin_allocated_WRITE_RD_0;
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port = FrontendPlugin_allocated_PHYS_RD_0;
  assign _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port = FrontendPlugin_allocated_ARCH_RD_0;
  assign _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port = FrontendPlugin_allocated_PHYS_RD_FREE_0;
  assign _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port = FrontendPlugin_allocated_BRANCH_SEL_0;
  assign _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port = FrontendPlugin_dispatch_Prediction_IS_BRANCH_0;
  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port_1 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_port = EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  assign _zz_RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_port_1 = (EU0_ExecutionUnitBase_pipeline_execute_1_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port = FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_0;
  assign _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port = FrontendPlugin_dispatch_LQ_ALLOC_0;
  assign _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_1 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port = FrontendPlugin_dispatch_SQ_ALLOC_0;
  assign _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_1 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port = FrontendPlugin_allocated_PHYS_RS_0_0;
  assign _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port = FrontendPlugin_allocated_READ_RS_0_0;
  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port = FrontendPlugin_allocated_PHYS_RS_1_0;
  assign _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port = FrontendPlugin_allocated_READ_RS_1_0;
  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port = FrontendPlugin_allocated_BRANCH_ID_0;
  assign _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port = FrontendPlugin_dispatch_LSU_ID_0;
  assign _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port_1 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port = FrontendPlugin_allocated_ROB_MSB_0;
  assign _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_AlignerPlugin_logic_extractors_0_pcWord_1 = AlignerPlugin_logic_extractors_0_firstWord;
  assign _zz_CommitDebugFilterPlugin_logic_commits_1 = CommitPlugin_logic_commit_event_mask[0];
  assign _zz_BranchContextPlugin_logic_onCommit_commitedNext_2 = BranchContextPlugin_logic_onCommit_isBranchCommit_0;
  assign _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount_1 = Lsu2Plugin_logic_lq_onCommit_lqCommits_0;
  assign _zz_Lsu2Plugin_logic_allocation_loads_requestsCount_1 = Lsu2Plugin_logic_allocation_loads_requests_0;
  assign _zz_Lsu2Plugin_logic_allocation_stores_requestsCount_1 = Lsu2Plugin_logic_allocation_stores_requests_0;
  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_1 = Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress[1 : 0];
  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_3 = Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress[1 : 1];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits = (! Lsu2Plugin_setup_specialTrap_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_1 = (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_1_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_2 = (! CommitPlugin_logic_reschedule_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_3 = (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age < CommitPlugin_logic_reschedule_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_4 = (! Lsu2Plugin_setup_sharedTrap_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_5 = (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_6 = (! CommitPlugin_logic_reschedule_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_7 = (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age < CommitPlugin_logic_reschedule_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_8 = (! Lsu2Plugin_setup_sharedTrap_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_9 = (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_10 = (! CommitPlugin_logic_reschedule_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_11 = (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age < CommitPlugin_logic_reschedule_age);
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_1 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[9];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_2 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[10];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_3 = {ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[11],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[12],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[13],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[14],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[15],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[16],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[17],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[18],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[19],{_zz_ALU0_ShiftPlugin_logic_process_reversed_4,{_zz_ALU0_ShiftPlugin_logic_process_reversed_5,_zz_ALU0_ShiftPlugin_logic_process_reversed_6}}}}}}}}}}};
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_4 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[20];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_5 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[21];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_6 = {ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[22],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[23],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[24],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[25],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[26],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[27],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[28],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[29],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[30],ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]}}}}}}}}};
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_1 = ALU0_ShiftPlugin_logic_process_shifted[9];
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_2 = ALU0_ShiftPlugin_logic_process_shifted[10];
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_3 = {ALU0_ShiftPlugin_logic_process_shifted[11],{ALU0_ShiftPlugin_logic_process_shifted[12],{ALU0_ShiftPlugin_logic_process_shifted[13],{ALU0_ShiftPlugin_logic_process_shifted[14],{ALU0_ShiftPlugin_logic_process_shifted[15],{ALU0_ShiftPlugin_logic_process_shifted[16],{ALU0_ShiftPlugin_logic_process_shifted[17],{ALU0_ShiftPlugin_logic_process_shifted[18],{ALU0_ShiftPlugin_logic_process_shifted[19],{_zz_ALU0_ShiftPlugin_logic_process_patched_4,{_zz_ALU0_ShiftPlugin_logic_process_patched_5,_zz_ALU0_ShiftPlugin_logic_process_patched_6}}}}}}}}}}};
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_4 = ALU0_ShiftPlugin_logic_process_shifted[20];
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_5 = ALU0_ShiftPlugin_logic_process_shifted[21];
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_6 = {ALU0_ShiftPlugin_logic_process_shifted[22],{ALU0_ShiftPlugin_logic_process_shifted[23],{ALU0_ShiftPlugin_logic_process_shifted[24],{ALU0_ShiftPlugin_logic_process_shifted[25],{ALU0_ShiftPlugin_logic_process_shifted[26],{ALU0_ShiftPlugin_logic_process_shifted[27],{ALU0_ShiftPlugin_logic_process_shifted[28],{ALU0_ShiftPlugin_logic_process_shifted[29],{ALU0_ShiftPlugin_logic_process_shifted[30],ALU0_ShiftPlugin_logic_process_shifted[31]}}}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_1 = 3'b010;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_2 = (3'b001 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_3 = (3'b000 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_1 = 3'b010;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_2 = (3'b001 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_3 = (3'b000 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_1 = 3'b010;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_2 = (3'b001 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_3 = (3'b000 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_1 = 3'b010;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_2 = (3'b001 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_3 = (3'b000 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_physicalAddress,_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_1};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_2 = 32'h00000000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_3 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_physicalAddress,_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_4};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_5 = 32'h00000000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_6 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_physicalAddress,_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_7};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_8 = 32'h00000000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_9 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_physicalAddress,_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_10};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_11 = 32'h00000000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_12 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[21 : 0]};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_13 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[21 : 0]};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_1 = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_4 = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_7 = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_10 = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0];
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented = COMB_CSR_770;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_1 = {COMB_CSR_772,{COMB_CSR_836,{COMB_CSR_768,{COMB_CSR_834,{COMB_CSR_769,{COMB_CSR_3860,{COMB_CSR_3859,{COMB_CSR_3858,{COMB_CSR_3857,{COMB_CSR_832,{_zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_2,_zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_3}}}}}}}}}}};
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_2 = COMB_CSR_833;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_3 = {COMB_CSR_835,COMB_CSR_773};
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated = {FetchPlugin_stages_1_MMU_L0_ENTRIES_0_physicalAddress,_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_1};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_2 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_3 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_1_physicalAddress,_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_4};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_5 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_6 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_2_physicalAddress,_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_7};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_8 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_9 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_3_physicalAddress,_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_10};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_11 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_12 = {FetchPlugin_stages_1_MMU_L1_ENTRIES_0_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[21 : 0]};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_13 = {FetchPlugin_stages_1_MMU_L1_ENTRIES_1_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[21 : 0]};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_1 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_4 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_7 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_10 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0];
  assign _zz_FrontendPlugin_decoded_LEGAL_0 = 32'h0000107f;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_1 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000207f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_2 = 32'h00002073;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_3 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000407f) == 32'h00004063);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_4 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000207f) == 32'h00002013);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_5 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000107f) == 32'h00000013),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000603f) == 32'h00000023),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_LEGAL_0_6) == 32'h00000003),{(_zz_FrontendPlugin_decoded_LEGAL_0_7 == _zz_FrontendPlugin_decoded_LEGAL_0_8),{_zz_FrontendPlugin_decoded_LEGAL_0_9,{_zz_FrontendPlugin_decoded_LEGAL_0_10,_zz_FrontendPlugin_decoded_LEGAL_0_11}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_0_6 = 32'h0000207f;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_7 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000505f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_8 = 32'h00000003;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_9 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000707b) == 32'h00000063);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_10 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000607f) == 32'h0000000f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_11 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h1800707f) == 32'h0000202f),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hfc00007f) == 32'h00000033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_LEGAL_0_12) == 32'h0800202f),{(_zz_FrontendPlugin_decoded_LEGAL_0_13 == _zz_FrontendPlugin_decoded_LEGAL_0_14),{_zz_FrontendPlugin_decoded_LEGAL_0_15,{_zz_FrontendPlugin_decoded_LEGAL_0_16,_zz_FrontendPlugin_decoded_LEGAL_0_17}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_0_12 = 32'he800707f;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_13 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hfc00305f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_14 = 32'h00001013;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_15 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h01f0707f) == 32'h0000500f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_16 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hbc00707f) == 32'h00005013);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_17 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hbe00707f) == 32'h00005033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hbe00707f) == 32'h00000033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_LEGAL_0_18) == 32'h1000202f),{(_zz_FrontendPlugin_decoded_LEGAL_0_19 == _zz_FrontendPlugin_decoded_LEGAL_0_20),{_zz_FrontendPlugin_decoded_LEGAL_0_21,{_zz_FrontendPlugin_decoded_LEGAL_0_22,_zz_FrontendPlugin_decoded_LEGAL_0_23}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_0_18 = 32'hf9f0707f;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_19 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hfe007fff);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_20 = 32'h12000073;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_21 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hdfffffff) == 32'h10200073);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_22 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hffefffff) == 32'h00000073);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_23 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hffffffff) == 32'h10500073);
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_2 = 32'h00002008;
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_3 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000050);
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_4 = 32'h00000010;
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_5 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000000c) == 32'h00000004);
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_6 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000028) == 32'h00000000);
  always @(posedge clk) begin
    if(_zz_30) begin
      FetchCachePlugin_logic_banks_0_mem[FetchCachePlugin_logic_banks_0_write_payload_address] <= FetchCachePlugin_logic_banks_0_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchCachePlugin_logic_banks_0_read_cmd_valid) begin
      FetchCachePlugin_logic_banks_0_mem_spinal_port1 <= FetchCachePlugin_logic_banks_0_mem[FetchCachePlugin_logic_banks_0_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_logic_ways_0_mem_port_1) begin
      FetchCachePlugin_logic_ways_0_mem[FetchCachePlugin_logic_waysWrite_address] <= _zz_FetchCachePlugin_logic_ways_0_mem_port;
    end
  end

  assign FetchCachePlugin_logic_ways_0_mem_spinal_port1 = FetchCachePlugin_logic_ways_0_mem[FetchCachePlugin_logic_ways_0_read_cmd_payload];
  always @(posedge clk) begin
    if(_zz_29) begin
      BranchContextPlugin_logic_mem_earlyBranch[FrontendPlugin_allocated_BRANCH_ID_0] <= _zz_BranchContextPlugin_logic_mem_earlyBranch_port;
    end
  end

  assign BranchContextPlugin_logic_mem_earlyBranch_spinal_port1 = BranchContextPlugin_logic_mem_earlyBranch[EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID];
  always @(posedge clk) begin
    if(_zz_8) begin
      BranchContextPlugin_logic_mem_finalBranch[EU0_BranchPlugin_logic_branch_finalBranch_payload_address] <= _zz_BranchContextPlugin_logic_mem_finalBranch_port;
    end
  end

  assign BranchContextPlugin_logic_mem_finalBranch_spinal_port1 = BranchContextPlugin_logic_mem_finalBranch[BranchContextPlugin_free_learn_bid];
  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_DecoderPredictionPlugin_logic_ras_mem_stack.bin",DecoderPredictionPlugin_logic_ras_mem_stack);
  end
  assign DecoderPredictionPlugin_logic_ras_mem_stack_spinal_port0 = DecoderPredictionPlugin_logic_ras_mem_stack[DecoderPredictionPlugin_logic_ras_ptr_pop];
  always @(posedge clk) begin
    if(_zz_28) begin
      DecoderPredictionPlugin_logic_ras_mem_stack[DecoderPredictionPlugin_logic_ras_write_payload_address] <= _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port;
    end
  end

  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_BtbPlugin_logic_mem.bin",BtbPlugin_logic_mem);
  end
  always @(posedge clk) begin
    if(FetchPlugin_stages_0_ready) begin
      BtbPlugin_logic_mem_spinal_port1 <= BtbPlugin_logic_mem[BtbPlugin_logic_readCmd_entryAddress];
    end
    if(_zz_27) begin
      BtbPlugin_logic_mem[BtbPlugin_logic_onLearn_port_payload_address] <= _zz_BtbPlugin_logic_mem_port;
    end
  end

  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_GSharePlugin_logic_mem_counter.bin",GSharePlugin_logic_mem_counter);
  end
  always @(posedge clk) begin
    if(_zz_26) begin
      GSharePlugin_logic_mem_counter[GSharePlugin_logic_mem_write_payload_address] <= _zz_GSharePlugin_logic_mem_counter_port;
    end
  end

  always @(posedge clk) begin
    if(FetchPlugin_stages_0_ready) begin
      GSharePlugin_logic_mem_counter_spinal_port1 <= GSharePlugin_logic_mem_counter[FetchPlugin_stages_0_GSharePlugin_logic_HASH];
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_addressPre[_zz_Lsu2Plugin_logic_lq_mem_addressPre_port] <= _zz_Lsu2Plugin_logic_lq_mem_addressPre_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_addressPre_spinal_port1 = Lsu2Plugin_logic_lq_mem_addressPre[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign Lsu2Plugin_logic_lq_mem_addressPre_spinal_port2 = Lsu2Plugin_logic_lq_mem_addressPre[Lsu2Plugin_logic_lq_ptr_freeReal];
  assign Lsu2Plugin_logic_lq_mem_addressPost_spinal_port0 = Lsu2Plugin_logic_lq_mem_addressPost[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(_zz_16) begin
      Lsu2Plugin_logic_lq_mem_addressPost[Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID] <= _zz_Lsu2Plugin_logic_lq_mem_addressPost_port;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_addressPost_spinal_port2 = Lsu2Plugin_logic_lq_mem_addressPost[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_size[_zz_Lsu2Plugin_logic_lq_mem_size_port] <= _zz_Lsu2Plugin_logic_lq_mem_size_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_size_spinal_port1 = Lsu2Plugin_logic_lq_mem_size[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign Lsu2Plugin_logic_lq_mem_size_spinal_port2 = Lsu2Plugin_logic_lq_mem_size[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_physRd[_zz_Lsu2Plugin_logic_lq_mem_physRd_port] <= _zz_Lsu2Plugin_logic_lq_mem_physRd_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_physRd_spinal_port1 = Lsu2Plugin_logic_lq_mem_physRd[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign Lsu2Plugin_logic_lq_mem_physRd_spinal_port2 = Lsu2Plugin_logic_lq_mem_physRd[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_robId[_zz_Lsu2Plugin_logic_lq_mem_robId_port] <= _zz_Lsu2Plugin_logic_lq_mem_robId_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_robId_spinal_port1 = Lsu2Plugin_logic_lq_mem_robId[Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID];
  assign Lsu2Plugin_logic_lq_mem_robId_spinal_port2 = Lsu2Plugin_logic_lq_mem_robId[Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel];
  assign Lsu2Plugin_logic_lq_mem_robId_spinal_port3 = Lsu2Plugin_logic_lq_mem_robId[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_robIdMsb[_zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port] <= _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_robIdMsb_spinal_port1 = Lsu2Plugin_logic_lq_mem_robIdMsb[Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_pc[_zz_Lsu2Plugin_logic_lq_mem_pc_port] <= _zz_Lsu2Plugin_logic_lq_mem_pc_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_pc_spinal_port1 = Lsu2Plugin_logic_lq_mem_pc[_zz_Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC];
  always @(posedge clk) begin
    if(_zz_23) begin
      Lsu2Plugin_logic_lq_mem_sqAlloc[FrontendPlugin_dispatch_LQ_ID_0] <= _zz_Lsu2Plugin_logic_lq_mem_sqAlloc_port;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port1 = Lsu2Plugin_logic_lq_mem_sqAlloc[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port2 = Lsu2Plugin_logic_lq_mem_sqAlloc[_zz_Lsu2Plugin_logic_lq_mem_sqAlloc_port_1];
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port3 = Lsu2Plugin_logic_lq_mem_sqAlloc[Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID];
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port4 = Lsu2Plugin_logic_lq_mem_sqAlloc[Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ID];
  assign Lsu2Plugin_logic_lq_mem_io_spinal_port0 = Lsu2Plugin_logic_lq_mem_io[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(_zz_15) begin
      Lsu2Plugin_logic_lq_mem_io[Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID] <= _zz_Lsu2Plugin_logic_lq_mem_io_port;
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_writeRd[_zz_Lsu2Plugin_logic_lq_mem_writeRd_port] <= _zz_Lsu2Plugin_logic_lq_mem_writeRd_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_writeRd_spinal_port1 = Lsu2Plugin_logic_lq_mem_writeRd[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign Lsu2Plugin_logic_lq_mem_writeRd_spinal_port2 = Lsu2Plugin_logic_lq_mem_writeRd[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_lr[_zz_Lsu2Plugin_logic_lq_mem_lr_port] <= _zz_Lsu2Plugin_logic_lq_mem_lr_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_lr_spinal_port1 = Lsu2Plugin_logic_lq_mem_lr[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_unsigned[_zz_Lsu2Plugin_logic_lq_mem_unsigned_port] <= _zz_Lsu2Plugin_logic_lq_mem_unsigned_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_unsigned_spinal_port1 = Lsu2Plugin_logic_lq_mem_unsigned[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign Lsu2Plugin_logic_lq_mem_unsigned_spinal_port2 = Lsu2Plugin_logic_lq_mem_unsigned[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(_zz_22) begin
      Lsu2Plugin_logic_lq_mem_doSpecial[FrontendPlugin_dispatch_LQ_ID_0] <= _zz_Lsu2Plugin_logic_lq_mem_doSpecial_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_10) begin
      Lsu2Plugin_logic_lq_mem_doSpecial[Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID] <= _zz_Lsu2Plugin_logic_lq_mem_doSpecial_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_doSpecial_spinal_port2 = Lsu2Plugin_logic_lq_mem_doSpecial[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_needTranslation[_zz_Lsu2Plugin_logic_lq_mem_needTranslation_port] <= _zz_Lsu2Plugin_logic_lq_mem_needTranslation_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_needTranslation_spinal_port1 = Lsu2Plugin_logic_lq_mem_needTranslation[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(_zz_14) begin
      Lsu2Plugin_logic_lq_mem_needTranslation[Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID] <= _zz_Lsu2Plugin_logic_lq_mem_needTranslation_port_2;
    end
  end

  always @(posedge clk) begin
    if(_zz_21) begin
      Lsu2Plugin_logic_lq_mem_spFpAddress[FrontendPlugin_dispatch_LQ_ID_0] <= _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port;
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_hazardPrediction_valid[_zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port] <= _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_spinal_port1 = Lsu2Plugin_logic_lq_mem_hazardPrediction_valid[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_hazardPrediction_delta[_zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port] <= _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_spinal_port1 = Lsu2Plugin_logic_lq_mem_hazardPrediction_delta[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_hazardPrediction_score[_zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port] <= _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port_1;
    end
  end

  assign Lsu2Plugin_logic_lq_mem_hazardPrediction_score_spinal_port1 = Lsu2Plugin_logic_lq_mem_hazardPrediction_score[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_hitPrediction_counter[_zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port] <= _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port_1;
    end
  end

  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_Lsu2Plugin_logic_lq_hazardPrediction_mem.bin",Lsu2Plugin_logic_lq_hazardPrediction_mem);
  end
  always @(posedge clk) begin
    if(_zz_25) begin
      Lsu2Plugin_logic_lq_hazardPrediction_mem[Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_address] <= _zz_Lsu2Plugin_logic_lq_hazardPrediction_mem_port;
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_valid) begin
      Lsu2Plugin_logic_lq_hazardPrediction_mem_spinal_port1 <= Lsu2Plugin_logic_lq_hazardPrediction_mem[Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_payload];
    end
  end

  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_Lsu2Plugin_logic_lq_hitPrediction_mem.bin",Lsu2Plugin_logic_lq_hitPrediction_mem);
  end
  always @(posedge clk) begin
    if(_zz_24) begin
      Lsu2Plugin_logic_lq_hitPrediction_mem[Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_address] <= _zz_Lsu2Plugin_logic_lq_hitPrediction_mem_port;
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_valid) begin
      Lsu2Plugin_logic_lq_hitPrediction_mem_spinal_port1 <= Lsu2Plugin_logic_lq_hitPrediction_mem[Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_robId[_zz_Lsu2Plugin_logic_sq_mem_robId_port] <= _zz_Lsu2Plugin_logic_sq_mem_robId_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_robId_spinal_port1 = Lsu2Plugin_logic_sq_mem_robId[Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID];
  assign Lsu2Plugin_logic_sq_mem_robId_spinal_port2 = Lsu2Plugin_logic_sq_mem_robId[Lsu2Plugin_logic_sq_ptr_commitReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_robIdMsb[_zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port] <= _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_robIdMsb_spinal_port1 = Lsu2Plugin_logic_sq_mem_robIdMsb[Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_addressPre[_zz_Lsu2Plugin_logic_sq_mem_addressPre_port] <= _zz_Lsu2Plugin_logic_sq_mem_addressPre_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_addressPre_spinal_port1 = Lsu2Plugin_logic_sq_mem_addressPre[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  assign Lsu2Plugin_logic_sq_mem_addressPre_spinal_port2 = Lsu2Plugin_logic_sq_mem_addressPre[Lsu2Plugin_logic_sq_ptr_commitReal];
  assign Lsu2Plugin_logic_sq_mem_addressPost_spinal_port0 = Lsu2Plugin_logic_sq_mem_addressPost[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  always @(posedge clk) begin
    if(_zz_13) begin
      Lsu2Plugin_logic_sq_mem_addressPost[Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID] <= _zz_Lsu2Plugin_logic_sq_mem_addressPost_port;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_addressPost_spinal_port2 = Lsu2Plugin_logic_sq_mem_addressPost[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  assign Lsu2Plugin_logic_sq_mem_addressPost_spinal_port3 = Lsu2Plugin_logic_sq_mem_addressPost[Lsu2Plugin_logic_sq_ptr_writeBackReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_size[_zz_Lsu2Plugin_logic_sq_mem_size_port] <= _zz_Lsu2Plugin_logic_sq_mem_size_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_size_spinal_port1 = Lsu2Plugin_logic_sq_mem_size[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  assign Lsu2Plugin_logic_sq_mem_size_spinal_port2 = Lsu2Plugin_logic_sq_mem_size[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  assign Lsu2Plugin_logic_sq_mem_size_spinal_port3 = Lsu2Plugin_logic_sq_mem_size[Lsu2Plugin_logic_sq_ptr_writeBackReal];
  assign Lsu2Plugin_logic_sq_mem_size_spinal_port4 = Lsu2Plugin_logic_sq_mem_size[Lsu2Plugin_logic_sq_ptr_commitReal];
  assign Lsu2Plugin_logic_sq_mem_io_spinal_port0 = Lsu2Plugin_logic_sq_mem_io[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  always @(posedge clk) begin
    if(_zz_12) begin
      Lsu2Plugin_logic_sq_mem_io[Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID] <= _zz_Lsu2Plugin_logic_sq_mem_io_port;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_io_spinal_port2 = Lsu2Plugin_logic_sq_mem_io[Lsu2Plugin_logic_sq_ptr_writeBackReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_amo[_zz_Lsu2Plugin_logic_sq_mem_amo_port] <= _zz_Lsu2Plugin_logic_sq_mem_amo_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_amo_spinal_port1 = Lsu2Plugin_logic_sq_mem_amo[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  assign Lsu2Plugin_logic_sq_mem_amo_spinal_port2 = Lsu2Plugin_logic_sq_mem_amo[Lsu2Plugin_logic_sq_ptr_commitReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_sc[_zz_Lsu2Plugin_logic_sq_mem_sc_port] <= _zz_Lsu2Plugin_logic_sq_mem_sc_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_sc_spinal_port1 = Lsu2Plugin_logic_sq_mem_sc[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  assign Lsu2Plugin_logic_sq_mem_sc_spinal_port2 = Lsu2Plugin_logic_sq_mem_sc[Lsu2Plugin_logic_sq_ptr_commitReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_data[_zz_Lsu2Plugin_logic_sq_mem_data_port] <= AguPlugin_setup_port_payload_data;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_data_spinal_port1 = Lsu2Plugin_logic_sq_mem_data[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  assign Lsu2Plugin_logic_sq_mem_data_spinal_port2 = Lsu2Plugin_logic_sq_mem_data[Lsu2Plugin_logic_sq_ptr_writeBackReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_needTranslation[_zz_Lsu2Plugin_logic_sq_mem_needTranslation_port] <= _zz_Lsu2Plugin_logic_sq_mem_needTranslation_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_needTranslation_spinal_port1 = Lsu2Plugin_logic_sq_mem_needTranslation[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  always @(posedge clk) begin
    if(_zz_11) begin
      Lsu2Plugin_logic_sq_mem_needTranslation[Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID] <= _zz_Lsu2Plugin_logic_sq_mem_needTranslation_port_2;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_needTranslation_spinal_port3 = Lsu2Plugin_logic_sq_mem_needTranslation[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  always @(posedge clk) begin
    if(_zz_18) begin
      Lsu2Plugin_logic_sq_mem_feededOnce[FrontendPlugin_dispatch_SQ_ID_0] <= _zz_Lsu2Plugin_logic_sq_mem_feededOnce_port;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_feededOnce_spinal_port1 = Lsu2Plugin_logic_sq_mem_feededOnce[Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SQID];
  always @(posedge clk) begin
    if(_zz_17) begin
      Lsu2Plugin_logic_sq_mem_feededOnce[Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID] <= _zz_Lsu2Plugin_logic_sq_mem_feededOnce_port_1;
    end
  end

  always @(posedge clk) begin
    if(_zz_20) begin
      Lsu2Plugin_logic_sq_mem_doSpecial[FrontendPlugin_dispatch_SQ_ID_0] <= _zz_Lsu2Plugin_logic_sq_mem_doSpecial_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_9) begin
      Lsu2Plugin_logic_sq_mem_doSpecial[Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID] <= _zz_Lsu2Plugin_logic_sq_mem_doSpecial_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_doSpecial_spinal_port2 = Lsu2Plugin_logic_sq_mem_doSpecial[Lsu2Plugin_logic_sq_ptr_commitReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_doNotBypass[_zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port] <= _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port_1;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_doNotBypass_spinal_port1 = Lsu2Plugin_logic_sq_mem_doNotBypass[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  always @(posedge clk) begin
    if(_zz_19) begin
      Lsu2Plugin_logic_sq_mem_lqAlloc[FrontendPlugin_dispatch_SQ_ID_0] <= _zz_Lsu2Plugin_logic_sq_mem_lqAlloc_port;
    end
  end

  assign Lsu2Plugin_logic_sq_mem_lqAlloc_spinal_port1 = Lsu2Plugin_logic_sq_mem_lqAlloc[Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0[FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port;
    end
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_spinal_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0[FetchCachePlugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1[FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port;
    end
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_spinal_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1[FetchCachePlugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2[FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port;
    end
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_spinal_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2[FetchCachePlugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3[FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port;
    end
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_spinal_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3[FetchCachePlugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0[FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port;
    end
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_spinal_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0[FetchCachePlugin_logic_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1[FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port;
    end
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_spinal_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1[FetchCachePlugin_logic_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0[Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port;
    end
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_spinal_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1[Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port;
    end
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_spinal_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2[Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port;
    end
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_spinal_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3[Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port;
    end
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_spinal_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0[Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port;
    end
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_spinal_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1[Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port;
    end
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_spinal_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_7) begin
      CsrRamPlugin_logic_mem[CsrRamPlugin_logic_writeLogic_port_payload_address] <= CsrRamPlugin_logic_writeLogic_port_payload_data;
    end
  end

  assign CsrRamPlugin_logic_mem_spinal_port1 = CsrRamPlugin_logic_mem[CsrRamPlugin_logic_readLogic_port_address];
  always @(posedge clk) begin
    if(_zz_6) begin
      BranchContextPlugin_free_dispatchMem_mem[BranchContextPlugin_free_dispatchMem_writes_0_port_payload_address] <= BranchContextPlugin_free_dispatchMem_writes_0_port_payload_data;
    end
  end

  assign BranchContextPlugin_free_dispatchMem_mem_spinal_port1 = BranchContextPlugin_free_dispatchMem_mem[BranchContextPlugin_free_learn_bid];
  always @(posedge clk) begin
    if(_zz_5) begin
      RobPlugin_logic_completionMem_target[RobPlugin_logic_completionMem_targetWrite_payload_address] <= RobPlugin_logic_completionMem_targetWrite_payload_data;
    end
  end

  assign RobPlugin_logic_completionMem_target_spinal_port1 = RobPlugin_logic_completionMem_target[RobPlugin_logic_completionMem_reads_0_targetRead_address];
  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_RobPlugin_logic_completionMem_hits_0.bin",RobPlugin_logic_completionMem_hits_0);
  end
  assign RobPlugin_logic_completionMem_hits_0_spinal_port0 = RobPlugin_logic_completionMem_hits_0[RobPlugin_logic_completionMem_init_0_robId];
  assign RobPlugin_logic_completionMem_hits_0_spinal_port1 = RobPlugin_logic_completionMem_hits_0[Lsu2Plugin_setup_sharedCompletion_payload_id];
  always @(posedge clk) begin
    if(_zz_4) begin
      RobPlugin_logic_completionMem_hits_0[Lsu2Plugin_setup_sharedCompletion_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_0_port;
    end
  end

  assign RobPlugin_logic_completionMem_hits_0_spinal_port3 = RobPlugin_logic_completionMem_hits_0[_zz_CommitPlugin_setup_robLineMask_mask];
  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_RobPlugin_logic_completionMem_hits_1.bin",RobPlugin_logic_completionMem_hits_1);
  end
  assign RobPlugin_logic_completionMem_hits_1_spinal_port0 = RobPlugin_logic_completionMem_hits_1[RobPlugin_logic_completionMem_init_0_robId];
  assign RobPlugin_logic_completionMem_hits_1_spinal_port1 = RobPlugin_logic_completionMem_hits_1[Lsu2Plugin_setup_specialCompletion_payload_id];
  always @(posedge clk) begin
    if(_zz_3) begin
      RobPlugin_logic_completionMem_hits_1[Lsu2Plugin_setup_specialCompletion_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_1_port;
    end
  end

  assign RobPlugin_logic_completionMem_hits_1_spinal_port3 = RobPlugin_logic_completionMem_hits_1[_zz_CommitPlugin_setup_robLineMask_mask];
  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_RobPlugin_logic_completionMem_hits_2.bin",RobPlugin_logic_completionMem_hits_2);
  end
  assign RobPlugin_logic_completionMem_hits_2_spinal_port0 = RobPlugin_logic_completionMem_hits_2[RobPlugin_logic_completionMem_init_0_robId];
  assign RobPlugin_logic_completionMem_hits_2_spinal_port1 = RobPlugin_logic_completionMem_hits_2[ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id];
  always @(posedge clk) begin
    if(_zz_2) begin
      RobPlugin_logic_completionMem_hits_2[ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_2_port;
    end
  end

  assign RobPlugin_logic_completionMem_hits_2_spinal_port3 = RobPlugin_logic_completionMem_hits_2[_zz_CommitPlugin_setup_robLineMask_mask];
  initial begin
    $readmemb("NaxRiscvAxi4LinuxPlicClint.v_toplevel_RobPlugin_logic_completionMem_hits_3.bin",RobPlugin_logic_completionMem_hits_3);
  end
  assign RobPlugin_logic_completionMem_hits_3_spinal_port0 = RobPlugin_logic_completionMem_hits_3[RobPlugin_logic_completionMem_init_0_robId];
  assign RobPlugin_logic_completionMem_hits_3_spinal_port1 = RobPlugin_logic_completionMem_hits_3[EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id];
  always @(posedge clk) begin
    if(_zz_1) begin
      RobPlugin_logic_completionMem_hits_3[EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_3_port;
    end
  end

  assign RobPlugin_logic_completionMem_hits_3_spinal_port3 = RobPlugin_logic_completionMem_hits_3[_zz_CommitPlugin_setup_robLineMask_mask];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_1) begin
      RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_spinal_port1 = RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0[_zz_CommitPlugin_logic_commit_active];
  assign RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_spinal_port2 = RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0[_zz_integer_RfAllocationPlugin_logic_push_mask_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PC_banks_0_port_1) begin
      RobPlugin_logic_storage_PC_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_PC_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_PC_banks_0_spinal_port1 = RobPlugin_logic_storage_PC_banks_0[_zz_commit_pc_0];
  assign RobPlugin_logic_storage_PC_banks_0_spinal_port2 = RobPlugin_logic_storage_PC_banks_0[_zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc];
  assign RobPlugin_logic_storage_PC_banks_0_spinal_port3 = RobPlugin_logic_storage_PC_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC];
  assign RobPlugin_logic_storage_PC_banks_0_spinal_port4 = RobPlugin_logic_storage_PC_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port_1) begin
      RobPlugin_logic_storage_WRITE_RD_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port1 = RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0];
  assign RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port2 = RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_integer_RfAllocationPlugin_logic_push_writeRd_0];
  assign RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port3 = RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD];
  assign RobPlugin_logic_storage_WRITE_RD_banks_0_spinal_port4 = RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_1) begin
      RobPlugin_logic_storage_PHYS_RD_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_PHYS_RD_banks_0_spinal_port1 = RobPlugin_logic_storage_PHYS_RD_banks_0[_zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0];
  assign RobPlugin_logic_storage_PHYS_RD_banks_0_spinal_port2 = RobPlugin_logic_storage_PHYS_RD_banks_0[_zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_1) begin
      RobPlugin_logic_storage_ARCH_RD_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_ARCH_RD_banks_0_spinal_port1 = RobPlugin_logic_storage_ARCH_RD_banks_0[_zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_1) begin
      RobPlugin_logic_storage_PHYS_RD_FREE_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_spinal_port1 = RobPlugin_logic_storage_PHYS_RD_FREE_banks_0[_zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_1) begin
      RobPlugin_logic_storage_BRANCH_SEL_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_BRANCH_SEL_banks_0_spinal_port1 = RobPlugin_logic_storage_BRANCH_SEL_banks_0[_zz_BranchContextPlugin_logic_onCommit_isBranch_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port_1) begin
      RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0[FrontendPlugin_dispatch_ROB_ID] <= _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_spinal_port1 = RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0[_zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0];
  assign RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_spinal_port2 = RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0[_zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_port_1) begin
      RobPlugin_logic_storage_BRANCH_TAKEN_banks_0[EU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID] <= _zz_RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_spinal_port1 = RobPlugin_logic_storage_BRANCH_TAKEN_banks_0[_zz_HistoryPlugin_logic_onCommit_isTaken_0];
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_spinal_port2 = RobPlugin_logic_storage_BRANCH_TAKEN_banks_0[_zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port) begin
      RobPlugin_logic_storage_BRANCH_HISTORY_banks_0[FrontendPlugin_allocated_ROB_ID] <= FrontendPlugin_allocated_BRANCH_HISTORY_0;
    end
  end

  assign RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_spinal_port1 = RobPlugin_logic_storage_BRANCH_HISTORY_banks_0[_zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port_1) begin
      RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_spinal_port1 = RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0[_zz_DecoderPredictionPlugin_logic_ras_healPush];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_1) begin
      RobPlugin_logic_storage_LQ_ALLOC_banks_0[FrontendPlugin_dispatch_ROB_ID] <= _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_LQ_ALLOC_banks_0_spinal_port1 = RobPlugin_logic_storage_LQ_ALLOC_banks_0[_zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_1) begin
      RobPlugin_logic_storage_SQ_ALLOC_banks_0[FrontendPlugin_dispatch_ROB_ID] <= _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_SQ_ALLOC_banks_0_spinal_port1 = RobPlugin_logic_storage_SQ_ALLOC_banks_0[_zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port) begin
      RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0[FrontendPlugin_allocated_ROB_ID] <= FrontendPlugin_allocated_Frontend_MICRO_OP_0;
    end
  end

  assign RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_spinal_port1 = RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP];
  assign RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_spinal_port2 = RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port_1) begin
      RobPlugin_logic_storage_PHYS_RS_0_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_PHYS_RS_0_banks_0_spinal_port1 = RobPlugin_logic_storage_PHYS_RS_0_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port_1) begin
      RobPlugin_logic_storage_READ_RS_0_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_READ_RS_0_banks_0_spinal_port1 = RobPlugin_logic_storage_READ_RS_0_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0];
  assign RobPlugin_logic_storage_READ_RS_0_banks_0_spinal_port2 = RobPlugin_logic_storage_READ_RS_0_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port_1) begin
      RobPlugin_logic_storage_PHYS_RS_1_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_PHYS_RS_1_banks_0_spinal_port1 = RobPlugin_logic_storage_PHYS_RS_1_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port_1) begin
      RobPlugin_logic_storage_READ_RS_1_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_READ_RS_1_banks_0_spinal_port1 = RobPlugin_logic_storage_READ_RS_1_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1];
  assign RobPlugin_logic_storage_READ_RS_1_banks_0_spinal_port2 = RobPlugin_logic_storage_READ_RS_1_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port_1) begin
      RobPlugin_logic_storage_BRANCH_ID_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_BRANCH_ID_banks_0_spinal_port1 = RobPlugin_logic_storage_BRANCH_ID_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_LSU_ID_banks_0_port_1) begin
      RobPlugin_logic_storage_LSU_ID_banks_0[FrontendPlugin_dispatch_ROB_ID] <= _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_LSU_ID_banks_0_spinal_port1 = RobPlugin_logic_storage_LSU_ID_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port_1) begin
      RobPlugin_logic_storage_ROB_MSB_banks_0[FrontendPlugin_allocated_ROB_ID] <= _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port;
    end
  end

  assign RobPlugin_logic_storage_ROB_MSB_banks_0_spinal_port1 = RobPlugin_logic_storage_ROB_MSB_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB];
  AxiLite4Clint clintCtrl (
    .io_bus_aw_valid        (clint_awvalid                        ), //i
    .io_bus_aw_ready        (clintCtrl_io_bus_aw_ready            ), //o
    .io_bus_aw_payload_addr (clint_awaddr[15:0]                   ), //i
    .io_bus_aw_payload_prot (clint_awprot[2:0]                    ), //i
    .io_bus_w_valid         (clint_wvalid                         ), //i
    .io_bus_w_ready         (clintCtrl_io_bus_w_ready             ), //o
    .io_bus_w_payload_data  (clint_wdata[31:0]                    ), //i
    .io_bus_w_payload_strb  (clint_wstrb[3:0]                     ), //i
    .io_bus_b_valid         (clintCtrl_io_bus_b_valid             ), //o
    .io_bus_b_ready         (clint_bready                         ), //i
    .io_bus_b_payload_resp  (clintCtrl_io_bus_b_payload_resp[1:0] ), //o
    .io_bus_ar_valid        (clint_arvalid                        ), //i
    .io_bus_ar_ready        (clintCtrl_io_bus_ar_ready            ), //o
    .io_bus_ar_payload_addr (clint_araddr[15:0]                   ), //i
    .io_bus_ar_payload_prot (clint_arprot[2:0]                    ), //i
    .io_bus_r_valid         (clintCtrl_io_bus_r_valid             ), //o
    .io_bus_r_ready         (clint_rready                         ), //i
    .io_bus_r_payload_data  (clintCtrl_io_bus_r_payload_data[31:0]), //o
    .io_bus_r_payload_resp  (clintCtrl_io_bus_r_payload_resp[1:0] ), //o
    .io_timerInterrupt      (clintCtrl_io_timerInterrupt          ), //o
    .io_softwareInterrupt   (clintCtrl_io_softwareInterrupt       ), //o
    .io_time                (clintCtrl_io_time[63:0]              ), //o
    .clk                    (clk                                  ), //i
    .reset                  (reset                                )  //i
  );
  AxiLite4Plic plicCtrl (
    .io_bus_aw_valid        (plic_awvalid                        ), //i
    .io_bus_aw_ready        (plicCtrl_io_bus_aw_ready            ), //o
    .io_bus_aw_payload_addr (plic_awaddr[21:0]                   ), //i
    .io_bus_aw_payload_prot (plic_awprot[2:0]                    ), //i
    .io_bus_w_valid         (plic_wvalid                         ), //i
    .io_bus_w_ready         (plicCtrl_io_bus_w_ready             ), //o
    .io_bus_w_payload_data  (plic_wdata[31:0]                    ), //i
    .io_bus_w_payload_strb  (plic_wstrb[3:0]                     ), //i
    .io_bus_b_valid         (plicCtrl_io_bus_b_valid             ), //o
    .io_bus_b_ready         (plic_bready                         ), //i
    .io_bus_b_payload_resp  (plicCtrl_io_bus_b_payload_resp[1:0] ), //o
    .io_bus_ar_valid        (plic_arvalid                        ), //i
    .io_bus_ar_ready        (plicCtrl_io_bus_ar_ready            ), //o
    .io_bus_ar_payload_addr (plic_araddr[21:0]                   ), //i
    .io_bus_ar_payload_prot (plic_arprot[2:0]                    ), //i
    .io_bus_r_valid         (plicCtrl_io_bus_r_valid             ), //o
    .io_bus_r_ready         (plic_rready                         ), //i
    .io_bus_r_payload_data  (plicCtrl_io_bus_r_payload_data[31:0]), //o
    .io_bus_r_payload_resp  (plicCtrl_io_bus_r_payload_resp[1:0] ), //o
    .io_sources             (plicCtrl_io_sources[30:0]           ), //i
    .io_targets             (plicCtrl_io_targets[1:0]            ), //o
    .clk                    (clk                                 ), //i
    .reset                  (reset                               )  //i
  );
  TranslatorWithRollback integer_RfTranslationPlugin_logic_impl (
    .io_rollback                  (integer_RfTranslationPlugin_logic_impl_io_rollback                      ), //i
    .io_writes_0_valid            (integer_RfTranslationPlugin_logic_impl_io_writes_0_valid                ), //i
    .io_writes_0_payload_address  (FrontendPlugin_allocated_ARCH_RD_0[4:0]                                 ), //i
    .io_writes_0_payload_data     (FrontendPlugin_allocated_PHYS_RD_0[5:0]                                 ), //i
    .io_commits_0_valid           (integer_RfTranslationPlugin_logic_impl_io_commits_0_valid               ), //i
    .io_commits_0_payload_address (integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_address[4:0]), //i
    .io_commits_0_payload_data    (integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_data[5:0]   ), //i
    .io_reads_0_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_0_cmd_valid             ), //i
    .io_reads_0_cmd_payload       (FrontendPlugin_allocated_ARCH_RD_0[4:0]                                 ), //i
    .io_reads_0_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_valid             ), //o
    .io_reads_0_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_payload[5:0]      ), //o
    .io_reads_1_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_1_cmd_valid             ), //i
    .io_reads_1_cmd_payload       (FrontendPlugin_allocated_ARCH_RS_0_0[4:0]                               ), //i
    .io_reads_1_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_valid             ), //o
    .io_reads_1_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_payload[5:0]      ), //o
    .io_reads_2_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_2_cmd_valid             ), //i
    .io_reads_2_cmd_payload       (FrontendPlugin_allocated_ARCH_RS_1_0[4:0]                               ), //i
    .io_reads_2_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_valid             ), //o
    .io_reads_2_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_payload[5:0]      ), //o
    .clk                          (clk                                                                     ), //i
    .reset                        (reset                                                                   )  //i
  );
  AllocatorMultiPortMem integer_RfAllocationPlugin_logic_allocator (
    .io_push_0_valid   (integer_RfAllocationPlugin_logic_allocator_io_push_0_valid       ), //i
    .io_push_0_payload (integer_RfAllocationPlugin_logic_allocator_io_push_0_payload[5:0]), //i
    .io_pop_mask       (integer_RfAllocationPlugin_logic_allocator_io_pop_mask           ), //i
    .io_pop_ready      (integer_RfAllocationPlugin_logic_allocator_io_pop_ready          ), //o
    .io_pop_fire       (FrontendPlugin_allocated_isFireing                               ), //i
    .io_pop_values_0   (integer_RfAllocationPlugin_logic_allocator_io_pop_values_0[5:0]  ), //o
    .clk               (clk                                                              ), //i
    .reset             (reset                                                            )  //i
  );
  DataCache DataCachePlugin_logic_cache (
    .io_lock_valid                             (DataCachePlugin_setup_lockPort_valid                                       ), //i
    .io_lock_address                           (DataCachePlugin_setup_lockPort_address[31:0]                               ), //i
    .io_load_cmd_valid                         (DataCachePlugin_logic_load_hit                                             ), //i
    .io_load_cmd_ready                         (DataCachePlugin_logic_cache_io_load_cmd_ready                              ), //o
    .io_load_cmd_payload_virtual               (DataCachePlugin_logic_cache_io_load_cmd_payload_virtual[31:0]              ), //i
    .io_load_cmd_payload_size                  (DataCachePlugin_logic_cache_io_load_cmd_payload_size[1:0]                  ), //i
    .io_load_cmd_payload_redoOnDataHazard      (DataCachePlugin_logic_cache_io_load_cmd_payload_redoOnDataHazard           ), //i
    .io_load_cmd_payload_unlocked              (DataCachePlugin_logic_cache_io_load_cmd_payload_unlocked                   ), //i
    .io_load_cmd_payload_unique                (DataCachePlugin_logic_cache_io_load_cmd_payload_unique                     ), //i
    .io_load_translated_physical               (DataCachePlugin_logic_cache_io_load_translated_physical[31:0]              ), //i
    .io_load_translated_abord                  (DataCachePlugin_logic_cache_io_load_translated_abord                       ), //i
    .io_load_cancels                           (DataCachePlugin_logic_cache_io_load_cancels[2:0]                           ), //i
    .io_load_rsp_valid                         (DataCachePlugin_logic_cache_io_load_rsp_valid                              ), //o
    .io_load_rsp_payload_data                  (DataCachePlugin_logic_cache_io_load_rsp_payload_data[31:0]                 ), //o
    .io_load_rsp_payload_fault                 (DataCachePlugin_logic_cache_io_load_rsp_payload_fault                      ), //o
    .io_load_rsp_payload_redo                  (DataCachePlugin_logic_cache_io_load_rsp_payload_redo                       ), //o
    .io_load_rsp_payload_refillSlot            (DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlot[1:0]            ), //o
    .io_load_rsp_payload_refillSlotAny         (DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlotAny              ), //o
    .io_store_cmd_valid                        (Lsu2Plugin_setup_cacheStore_cmd_valid                                      ), //i
    .io_store_cmd_ready                        (DataCachePlugin_logic_cache_io_store_cmd_ready                             ), //o
    .io_store_cmd_payload_address              (Lsu2Plugin_setup_cacheStore_cmd_payload_address[31:0]                      ), //i
    .io_store_cmd_payload_data                 (Lsu2Plugin_setup_cacheStore_cmd_payload_data[31:0]                         ), //i
    .io_store_cmd_payload_mask                 (Lsu2Plugin_setup_cacheStore_cmd_payload_mask[3:0]                          ), //i
    .io_store_cmd_payload_generation           (Lsu2Plugin_setup_cacheStore_cmd_payload_generation                         ), //i
    .io_store_cmd_payload_io                   (Lsu2Plugin_setup_cacheStore_cmd_payload_io                                 ), //i
    .io_store_cmd_payload_flush                (Lsu2Plugin_setup_cacheStore_cmd_payload_flush                              ), //i
    .io_store_cmd_payload_flushFree            (Lsu2Plugin_setup_cacheStore_cmd_payload_flushFree                          ), //i
    .io_store_cmd_payload_prefetch             (Lsu2Plugin_setup_cacheStore_cmd_payload_prefetch                           ), //i
    .io_store_rsp_valid                        (DataCachePlugin_logic_cache_io_store_rsp_valid                             ), //o
    .io_store_rsp_payload_fault                (DataCachePlugin_logic_cache_io_store_rsp_payload_fault                     ), //o
    .io_store_rsp_payload_redo                 (DataCachePlugin_logic_cache_io_store_rsp_payload_redo                      ), //o
    .io_store_rsp_payload_refillSlot           (DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlot[1:0]           ), //o
    .io_store_rsp_payload_refillSlotAny        (DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlotAny             ), //o
    .io_store_rsp_payload_generationKo         (DataCachePlugin_logic_cache_io_store_rsp_payload_generationKo              ), //o
    .io_store_rsp_payload_flush                (DataCachePlugin_logic_cache_io_store_rsp_payload_flush                     ), //o
    .io_store_rsp_payload_prefetch             (DataCachePlugin_logic_cache_io_store_rsp_payload_prefetch                  ), //o
    .io_store_rsp_payload_address              (DataCachePlugin_logic_cache_io_store_rsp_payload_address[31:0]             ), //o
    .io_store_rsp_payload_io                   (DataCachePlugin_logic_cache_io_store_rsp_payload_io                        ), //o
    .io_mem_read_cmd_valid                     (DataCachePlugin_logic_cache_io_mem_read_cmd_valid                          ), //o
    .io_mem_read_cmd_ready                     (DataCachePlugin_mem_read_cmd_ready                                         ), //i
    .io_mem_read_cmd_payload_id                (DataCachePlugin_logic_cache_io_mem_read_cmd_payload_id                     ), //o
    .io_mem_read_cmd_payload_address           (DataCachePlugin_logic_cache_io_mem_read_cmd_payload_address[31:0]          ), //o
    .io_mem_read_rsp_valid                     (DataCachePlugin_mem_read_rsp_valid                                         ), //i
    .io_mem_read_rsp_ready                     (DataCachePlugin_logic_cache_io_mem_read_rsp_ready                          ), //o
    .io_mem_read_rsp_payload_id                (DataCachePlugin_mem_read_rsp_payload_id                                    ), //i
    .io_mem_read_rsp_payload_data              (DataCachePlugin_mem_read_rsp_payload_data[31:0]                            ), //i
    .io_mem_read_rsp_payload_error             (DataCachePlugin_mem_read_rsp_payload_error                                 ), //i
    .io_mem_write_cmd_valid                    (DataCachePlugin_logic_cache_io_mem_write_cmd_valid                         ), //o
    .io_mem_write_cmd_ready                    (DataCachePlugin_mem_write_cmd_ready                                        ), //i
    .io_mem_write_cmd_payload_last             (DataCachePlugin_logic_cache_io_mem_write_cmd_payload_last                  ), //o
    .io_mem_write_cmd_payload_fragment_address (DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_address[31:0]), //o
    .io_mem_write_cmd_payload_fragment_data    (DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_data[31:0]   ), //o
    .io_mem_write_cmd_payload_fragment_id      (DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_id           ), //o
    .io_mem_write_rsp_valid                    (DataCachePlugin_mem_write_rsp_valid                                        ), //i
    .io_mem_write_rsp_payload_error            (DataCachePlugin_mem_write_rsp_payload_error                                ), //i
    .io_mem_write_rsp_payload_id               (DataCachePlugin_mem_write_rsp_payload_id                                   ), //i
    .io_refillCompletions                      (DataCachePlugin_logic_cache_io_refillCompletions[1:0]                      ), //o
    .io_refillEvent                            (DataCachePlugin_logic_cache_io_refillEvent                                 ), //o
    .io_writebackEvent                         (DataCachePlugin_logic_cache_io_writebackEvent                              ), //o
    .io_writebackBusy                          (DataCachePlugin_logic_cache_io_writebackBusy                               ), //o
    .io_tagEvent                               (DataCachePlugin_logic_cache_io_tagEvent                                    ), //o
    .clk                                       (clk                                                                        ), //i
    .reset                                     (reset                                                                      )  //i
  );
  StreamFifoLowLatency CommitPlugin_logic_free_lineEventStream_fifo (
    .io_push_valid         (CommitPlugin_logic_free_lineEventStream_valid                         ), //i
    .io_push_ready         (CommitPlugin_logic_free_lineEventStream_fifo_io_push_ready            ), //o
    .io_push_payload_robId (CommitPlugin_logic_free_lineEventStream_payload_robId[3:0]            ), //i
    .io_push_payload_mask  (CommitPlugin_logic_free_lineEventStream_payload_mask                  ), //i
    .io_pop_valid          (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_valid             ), //o
    .io_pop_ready          (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_ready             ), //i
    .io_pop_payload_robId  (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_robId[3:0]), //o
    .io_pop_payload_mask   (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_mask      ), //o
    .io_flush              (CommitPlugin_logic_free_lineEventStream_fifo_io_flush                 ), //i
    .io_occupancy          (CommitPlugin_logic_free_lineEventStream_fifo_io_occupancy[4:0]        ), //o
    .io_availability       (CommitPlugin_logic_free_lineEventStream_fifo_io_availability[4:0]     ), //o
    .clk                   (clk                                                                   ), //i
    .reset                 (reset                                                                 )  //i
  );
  DivRadix4 EU0_DivPlugin_logic_div (
    .io_flush              (EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed                          ), //i
    .io_cmd_valid          (EU0_DivPlugin_logic_div_io_cmd_valid                                        ), //i
    .io_cmd_ready          (EU0_DivPlugin_logic_div_io_cmd_ready                                        ), //o
    .io_cmd_payload_a      (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED[31:0]), //i
    .io_cmd_payload_b      (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED[31:0]), //i
    .io_rsp_valid          (EU0_DivPlugin_logic_div_io_rsp_valid                                        ), //o
    .io_rsp_ready          (EU0_ExecutionUnitBase_pipeline_execute_1_ready                              ), //i
    .io_rsp_payload_result (EU0_DivPlugin_logic_div_io_rsp_payload_result[34:0]                         ), //o
    .io_rsp_payload_remain (EU0_DivPlugin_logic_div_io_rsp_payload_remain[32:0]                         ), //o
    .clk                   (clk                                                                         ), //i
    .reset                 (reset                                                                       )  //i
  );
  PrefetchPredictor Lsu2Plugin_logic_prefetch_predictor (
    .io_learn_valid            (Lsu2Plugin_logic_prefetch_predictor_io_learn_valid                 ), //i
    .io_learn_payload_physical (Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_address[31:0]     ), //i
    .io_learn_payload_allocate (Lsu2Plugin_logic_prefetch_predictor_io_learn_payload_allocate      ), //i
    .io_prediction_cmd_valid   (Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_valid        ), //o
    .io_prediction_cmd_ready   (Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready        ), //i
    .io_prediction_cmd_payload (Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_payload[31:0]), //o
    .io_prediction_rsp_valid   (Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_valid        ), //i
    .io_prediction_rsp_payload (Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_payload      )  //i
  );
  IssueQueue DispatchPlugin_logic_queue (
    .io_clear                                   (CommitPlugin_logic_commit_reschedulePort_valid                       ), //i
    .io_events                                  (DispatchPlugin_logic_wake_optReduce_reduced[7:0]                     ), //i
    .io_push_valid                              (FrontendPlugin_dispatch_isFireing                                    ), //i
    .io_push_ready                              (DispatchPlugin_logic_queue_io_push_ready                             ), //o
    .io_push_payload_slots_0_event              (DispatchPlugin_logic_queue_io_push_payload_slots_0_event[7:0]        ), //i
    .io_push_payload_slots_0_sel                (DispatchPlugin_logic_queue_io_push_payload_slots_0_sel[1:0]          ), //i
    .io_push_payload_slots_0_context_staticWake (DispatchPlugin_logic_queue_io_push_payload_slots_0_context_staticWake), //i
    .io_push_payload_slots_0_context_physRd     (FrontendPlugin_dispatch_PHYS_RD_0[5:0]                               ), //i
    .io_push_payload_slots_0_context_robId      (DispatchPlugin_logic_queue_io_push_payload_slots_0_context_robId[3:0]), //i
    .io_push_payload_slots_0_context_euCtx_0    (FrontendPlugin_dispatch_PHYS_RS_0_0[5:0]                             ), //i
    .io_push_payload_slots_0_context_euCtx_1    (FrontendPlugin_dispatch_PHYS_RS_1_0[5:0]                             ), //i
    .io_schedules_0_valid                       (DispatchPlugin_logic_queue_io_schedules_0_valid                      ), //o
    .io_schedules_0_ready                       (DispatchPlugin_logic_pop_0_stagesList_0_ready                        ), //i
    .io_schedules_0_payload_event               (DispatchPlugin_logic_queue_io_schedules_0_payload_event[7:0]         ), //o
    .io_schedules_1_valid                       (DispatchPlugin_logic_queue_io_schedules_1_valid                      ), //o
    .io_schedules_1_ready                       (DispatchPlugin_logic_pop_1_stagesList_0_ready                        ), //i
    .io_schedules_1_payload_event               (DispatchPlugin_logic_queue_io_schedules_1_payload_event[7:0]         ), //o
    .io_contexts_0_staticWake                   (DispatchPlugin_logic_queue_io_contexts_0_staticWake                  ), //o
    .io_contexts_0_physRd                       (DispatchPlugin_logic_queue_io_contexts_0_physRd[5:0]                 ), //o
    .io_contexts_0_robId                        (DispatchPlugin_logic_queue_io_contexts_0_robId[3:0]                  ), //o
    .io_contexts_0_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_0_euCtx_0[5:0]                ), //o
    .io_contexts_0_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_0_euCtx_1[5:0]                ), //o
    .io_contexts_1_staticWake                   (DispatchPlugin_logic_queue_io_contexts_1_staticWake                  ), //o
    .io_contexts_1_physRd                       (DispatchPlugin_logic_queue_io_contexts_1_physRd[5:0]                 ), //o
    .io_contexts_1_robId                        (DispatchPlugin_logic_queue_io_contexts_1_robId[3:0]                  ), //o
    .io_contexts_1_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_1_euCtx_0[5:0]                ), //o
    .io_contexts_1_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_1_euCtx_1[5:0]                ), //o
    .io_contexts_2_staticWake                   (DispatchPlugin_logic_queue_io_contexts_2_staticWake                  ), //o
    .io_contexts_2_physRd                       (DispatchPlugin_logic_queue_io_contexts_2_physRd[5:0]                 ), //o
    .io_contexts_2_robId                        (DispatchPlugin_logic_queue_io_contexts_2_robId[3:0]                  ), //o
    .io_contexts_2_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_2_euCtx_0[5:0]                ), //o
    .io_contexts_2_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_2_euCtx_1[5:0]                ), //o
    .io_contexts_3_staticWake                   (DispatchPlugin_logic_queue_io_contexts_3_staticWake                  ), //o
    .io_contexts_3_physRd                       (DispatchPlugin_logic_queue_io_contexts_3_physRd[5:0]                 ), //o
    .io_contexts_3_robId                        (DispatchPlugin_logic_queue_io_contexts_3_robId[3:0]                  ), //o
    .io_contexts_3_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_3_euCtx_0[5:0]                ), //o
    .io_contexts_3_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_3_euCtx_1[5:0]                ), //o
    .io_contexts_4_staticWake                   (DispatchPlugin_logic_queue_io_contexts_4_staticWake                  ), //o
    .io_contexts_4_physRd                       (DispatchPlugin_logic_queue_io_contexts_4_physRd[5:0]                 ), //o
    .io_contexts_4_robId                        (DispatchPlugin_logic_queue_io_contexts_4_robId[3:0]                  ), //o
    .io_contexts_4_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_4_euCtx_0[5:0]                ), //o
    .io_contexts_4_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_4_euCtx_1[5:0]                ), //o
    .io_contexts_5_staticWake                   (DispatchPlugin_logic_queue_io_contexts_5_staticWake                  ), //o
    .io_contexts_5_physRd                       (DispatchPlugin_logic_queue_io_contexts_5_physRd[5:0]                 ), //o
    .io_contexts_5_robId                        (DispatchPlugin_logic_queue_io_contexts_5_robId[3:0]                  ), //o
    .io_contexts_5_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_5_euCtx_0[5:0]                ), //o
    .io_contexts_5_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_5_euCtx_1[5:0]                ), //o
    .io_contexts_6_staticWake                   (DispatchPlugin_logic_queue_io_contexts_6_staticWake                  ), //o
    .io_contexts_6_physRd                       (DispatchPlugin_logic_queue_io_contexts_6_physRd[5:0]                 ), //o
    .io_contexts_6_robId                        (DispatchPlugin_logic_queue_io_contexts_6_robId[3:0]                  ), //o
    .io_contexts_6_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_6_euCtx_0[5:0]                ), //o
    .io_contexts_6_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_6_euCtx_1[5:0]                ), //o
    .io_contexts_7_staticWake                   (DispatchPlugin_logic_queue_io_contexts_7_staticWake                  ), //o
    .io_contexts_7_physRd                       (DispatchPlugin_logic_queue_io_contexts_7_physRd[5:0]                 ), //o
    .io_contexts_7_robId                        (DispatchPlugin_logic_queue_io_contexts_7_robId[3:0]                  ), //o
    .io_contexts_7_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_7_euCtx_0[5:0]                ), //o
    .io_contexts_7_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_7_euCtx_1[5:0]                ), //o
    .io_usage                                   (DispatchPlugin_logic_queue_io_usage[7:0]                             ), //o
    .clk                                        (clk                                                                  ), //i
    .reset                                      (reset                                                                )  //i
  );
  RegFileLatch integer_RegFilePlugin_logic_regfile_latches (
    .io_writes_0_valid   (integer_RegFilePlugin_logic_writeMerges_0_bus_valid              ), //i
    .io_writes_0_address (integer_RegFilePlugin_logic_writeMerges_0_bus_address[5:0]       ), //i
    .io_writes_0_data    (integer_RegFilePlugin_logic_writeMerges_0_bus_data[31:0]         ), //i
    .io_writes_0_robId   (integer_RegFilePlugin_logic_writeMerges_0_bus_robId[3:0]         ), //i
    .io_writes_1_valid   (integer_RegFilePlugin_logic_writeMerges_1_bus_valid              ), //i
    .io_writes_1_address (integer_RegFilePlugin_logic_writeMerges_1_bus_address[5:0]       ), //i
    .io_writes_1_data    (integer_RegFilePlugin_logic_writeMerges_1_bus_data[31:0]         ), //i
    .io_writes_1_robId   (integer_RegFilePlugin_logic_writeMerges_1_bus_robId[3:0]         ), //i
    .io_reads_0_valid    (ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid        ), //i
    .io_reads_0_address  (ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address[5:0] ), //i
    .io_reads_0_data     (integer_RegFilePlugin_logic_regfile_latches_io_reads_0_data[31:0]), //o
    .io_reads_1_valid    (ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid        ), //i
    .io_reads_1_address  (ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address[5:0] ), //i
    .io_reads_1_data     (integer_RegFilePlugin_logic_regfile_latches_io_reads_1_data[31:0]), //o
    .io_reads_2_valid    (EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid         ), //i
    .io_reads_2_address  (EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address[5:0]  ), //i
    .io_reads_2_data     (integer_RegFilePlugin_logic_regfile_latches_io_reads_2_data[31:0]), //o
    .io_reads_3_valid    (EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid         ), //i
    .io_reads_3_address  (EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address[5:0]  ), //i
    .io_reads_3_data     (integer_RegFilePlugin_logic_regfile_latches_io_reads_3_data[31:0]), //o
    .clk                 (clk                                                              ), //i
    .reset               (reset                                                            )  //i
  );
  DependencyStorage RfDependencyPlugin_logic_forRf_integer_impl (
    .io_writes_0_valid             (RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_valid                 ), //i
    .io_writes_0_payload_physical  (FrontendPlugin_dispatch_PHYS_RD_0[5:0]                                        ), //i
    .io_writes_0_payload_robId     (RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_payload_robId[3:0]    ), //i
    .io_commits_0_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_valid                ), //i
    .io_commits_0_payload_physical (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_payload_physical[5:0]), //i
    .io_commits_1_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_1_valid                ), //i
    .io_commits_1_payload_physical (Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_payload_physical[5:0]        ), //i
    .io_commits_2_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_2_valid                ), //i
    .io_commits_2_payload_physical (Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_payload_physical[5:0]                  ), //i
    .io_commits_3_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_3_valid                ), //i
    .io_commits_3_payload_physical (Lsu2Plugin_logic_special_wakeRf_payload_physical[5:0]                         ), //i
    .io_commits_4_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_4_valid                ), //i
    .io_commits_4_payload_physical (EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_payload_physical[5:0]        ), //i
    .io_reads_0_cmd_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_cmd_valid              ), //i
    .io_reads_0_cmd_payload        (FrontendPlugin_dispatch_PHYS_RS_0_0[5:0]                                      ), //i
    .io_reads_0_rsp_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_valid              ), //o
    .io_reads_0_rsp_payload_enable (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_enable     ), //o
    .io_reads_0_rsp_payload_rob    (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_rob[3:0]   ), //o
    .io_reads_1_cmd_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_cmd_valid              ), //i
    .io_reads_1_cmd_payload        (FrontendPlugin_dispatch_PHYS_RS_1_0[5:0]                                      ), //i
    .io_reads_1_rsp_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_valid              ), //o
    .io_reads_1_rsp_payload_enable (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_enable     ), //o
    .io_reads_1_rsp_payload_rob    (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_rob[3:0]   ), //o
    .clk                           (clk                                                                           ), //i
    .reset                         (reset                                                                         )  //i
  );
  always @(*) begin
    case(_zz_AlignerPlugin_logic_extractors_0_pcWord_1)
      1'b0 : _zz_AlignerPlugin_logic_extractors_0_pcWord = AlignerPlugin_logic_buffer_pc;
      default : _zz_AlignerPlugin_logic_extractors_0_pcWord = AlignerPlugin_setup_s2m_Fetch_FETCH_PC;
    endcase
  end

  always @(*) begin
    case(_zz_CommitDebugFilterPlugin_logic_commits_1)
      1'b0 : _zz_CommitDebugFilterPlugin_logic_commits = 1'b0;
      default : _zz_CommitDebugFilterPlugin_logic_commits = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_BranchContextPlugin_logic_onCommit_commitedNext_2)
      1'b0 : _zz_BranchContextPlugin_logic_onCommit_commitedNext_1 = 1'b0;
      default : _zz_BranchContextPlugin_logic_onCommit_commitedNext_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount_1)
      1'b0 : _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount = 1'b0;
      default : _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_allocation_loads_requestsCount_1)
      1'b0 : _zz_Lsu2Plugin_logic_allocation_loads_requestsCount = 1'b0;
      default : _zz_Lsu2Plugin_logic_allocation_loads_requestsCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_allocation_stores_requestsCount_1)
      1'b0 : _zz_Lsu2Plugin_logic_allocation_stores_requestsCount = 1'b0;
      default : _zz_Lsu2Plugin_logic_allocation_stores_requestsCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_1)
      2'b00 : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_0;
      2'b01 : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_1;
      2'b10 : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_2;
      default : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_3)
      1'b0 : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_2 = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_1;
      default : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_2 = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3;
    endcase
  end

  always @(*) begin
    case(Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID)
      3'b000 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_0_niceHazard;
      3'b001 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_1_niceHazard;
      3'b010 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_2_niceHazard;
      3'b011 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_3_niceHazard;
      3'b100 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_4_niceHazard;
      3'b101 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_5_niceHazard;
      3'b110 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_6_niceHazard;
      default : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_7_niceHazard;
    endcase
  end

  always @(*) begin
    case(CsrRamPlugin_logic_writeLogic_sel)
      2'b00 : begin
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_address = EU0_CsrAccessPlugin_logic_ramWritePort_address;
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_data = EU0_CsrAccessPlugin_logic_ramWritePort_data;
      end
      2'b01 : begin
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_address = PrivilegedPlugin_setup_ramWrite_address;
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_data = PrivilegedPlugin_setup_ramWrite_data;
      end
      default : begin
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_address = CsrRamPlugin_setup_initPort_address;
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_data = CsrRamPlugin_setup_initPort_data;
      end
    endcase
  end

  always @(*) begin
    case(CsrRamPlugin_logic_readLogic_sel)
      1'b0 : _zz_CsrRamPlugin_logic_readLogic_port_address = EU0_CsrAccessPlugin_logic_ramReadPort_address;
      default : _zz_CsrRamPlugin_logic_readLogic_port_address = PrivilegedPlugin_setup_ramRead_address;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
      Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "TRAP_ALIGN ";
      Lsu2Plugin_CTRL_ENUM_MMU_REDO : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "MMU_REDO   ";
      Lsu2Plugin_CTRL_ENUM_TRAP_MMU : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "TRAP_MMU   ";
      Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "LOAD_HAZARD";
      Lsu2Plugin_CTRL_ENUM_LOAD_MISS : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "LOAD_MISS  ";
      Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "LOAD_FAILED";
      Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "TRAP_ACCESS";
      Lsu2Plugin_CTRL_ENUM_SUCCESS : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "SUCCESS    ";
      default : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "???????????";
    endcase
  end
  always @(*) begin
    case(Lsu2Plugin_logic_sharedPip_stages_2_CTRL)
      Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "TRAP_ALIGN ";
      Lsu2Plugin_CTRL_ENUM_MMU_REDO : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "MMU_REDO   ";
      Lsu2Plugin_CTRL_ENUM_TRAP_MMU : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "TRAP_MMU   ";
      Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "LOAD_HAZARD";
      Lsu2Plugin_CTRL_ENUM_LOAD_MISS : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "LOAD_MISS  ";
      Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "LOAD_FAILED";
      Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "TRAP_ACCESS";
      Lsu2Plugin_CTRL_ENUM_SUCCESS : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "SUCCESS    ";
      default : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "???????????";
    endcase
  end
  always @(*) begin
    case(EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "BOOT ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "IDLE ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "READ ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "WRITE";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "DONE ";
      default : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(EU0_CsrAccessPlugin_logic_fsm_stateNext)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "BOOT ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "IDLE ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "READ ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "WRITE";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "DONE ";
      default : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_BOOT : EnvCallPlugin_logic_flushes_stateReg_string = "BOOT           ";
      EnvCallPlugin_logic_flushes_enumDef_IDLE : EnvCallPlugin_logic_flushes_stateReg_string = "IDLE           ";
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : EnvCallPlugin_logic_flushes_stateReg_string = "RESCHEDULE     ";
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : EnvCallPlugin_logic_flushes_stateReg_string = "VMA_FETCH_FLUSH";
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : EnvCallPlugin_logic_flushes_stateReg_string = "VMA_FETCH_WAIT ";
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : EnvCallPlugin_logic_flushes_stateReg_string = "LSU_FLUSH      ";
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : EnvCallPlugin_logic_flushes_stateReg_string = "WAIT_LSU       ";
      default : EnvCallPlugin_logic_flushes_stateReg_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(EnvCallPlugin_logic_flushes_stateNext)
      EnvCallPlugin_logic_flushes_enumDef_BOOT : EnvCallPlugin_logic_flushes_stateNext_string = "BOOT           ";
      EnvCallPlugin_logic_flushes_enumDef_IDLE : EnvCallPlugin_logic_flushes_stateNext_string = "IDLE           ";
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : EnvCallPlugin_logic_flushes_stateNext_string = "RESCHEDULE     ";
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : EnvCallPlugin_logic_flushes_stateNext_string = "VMA_FETCH_FLUSH";
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : EnvCallPlugin_logic_flushes_stateNext_string = "VMA_FETCH_WAIT ";
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : EnvCallPlugin_logic_flushes_stateNext_string = "LSU_FLUSH      ";
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : EnvCallPlugin_logic_flushes_stateNext_string = "WAIT_LSU       ";
      default : EnvCallPlugin_logic_flushes_stateNext_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(Lsu2Plugin_logic_special_atomic_stateReg)
      Lsu2Plugin_logic_special_atomic_enumDef_BOOT : Lsu2Plugin_logic_special_atomic_stateReg_string = "BOOT      ";
      Lsu2Plugin_logic_special_atomic_enumDef_IDLE : Lsu2Plugin_logic_special_atomic_stateReg_string = "IDLE      ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD : Lsu2Plugin_logic_special_atomic_stateReg_string = "LOAD_CMD  ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP : Lsu2Plugin_logic_special_atomic_stateReg_string = "LOAD_RSP  ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY : Lsu2Plugin_logic_special_atomic_stateReg_string = "LOCK_DELAY";
      Lsu2Plugin_logic_special_atomic_enumDef_ALU : Lsu2Plugin_logic_special_atomic_stateReg_string = "ALU       ";
      Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION : Lsu2Plugin_logic_special_atomic_stateReg_string = "COMPLETION";
      Lsu2Plugin_logic_special_atomic_enumDef_SYNC : Lsu2Plugin_logic_special_atomic_stateReg_string = "SYNC      ";
      Lsu2Plugin_logic_special_atomic_enumDef_TRAP : Lsu2Plugin_logic_special_atomic_stateReg_string = "TRAP      ";
      Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT : Lsu2Plugin_logic_special_atomic_stateReg_string = "TRAP_WAIT ";
      default : Lsu2Plugin_logic_special_atomic_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(Lsu2Plugin_logic_special_atomic_stateNext)
      Lsu2Plugin_logic_special_atomic_enumDef_BOOT : Lsu2Plugin_logic_special_atomic_stateNext_string = "BOOT      ";
      Lsu2Plugin_logic_special_atomic_enumDef_IDLE : Lsu2Plugin_logic_special_atomic_stateNext_string = "IDLE      ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD : Lsu2Plugin_logic_special_atomic_stateNext_string = "LOAD_CMD  ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP : Lsu2Plugin_logic_special_atomic_stateNext_string = "LOAD_RSP  ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY : Lsu2Plugin_logic_special_atomic_stateNext_string = "LOCK_DELAY";
      Lsu2Plugin_logic_special_atomic_enumDef_ALU : Lsu2Plugin_logic_special_atomic_stateNext_string = "ALU       ";
      Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION : Lsu2Plugin_logic_special_atomic_stateNext_string = "COMPLETION";
      Lsu2Plugin_logic_special_atomic_enumDef_SYNC : Lsu2Plugin_logic_special_atomic_stateNext_string = "SYNC      ";
      Lsu2Plugin_logic_special_atomic_enumDef_TRAP : Lsu2Plugin_logic_special_atomic_stateNext_string = "TRAP      ";
      Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT : Lsu2Plugin_logic_special_atomic_stateNext_string = "TRAP_WAIT ";
      default : Lsu2Plugin_logic_special_atomic_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_BOOT : MmuPlugin_logic_refill_stateReg_string = "BOOT ";
      MmuPlugin_logic_refill_enumDef_IDLE : MmuPlugin_logic_refill_stateReg_string = "IDLE ";
      MmuPlugin_logic_refill_enumDef_INIT : MmuPlugin_logic_refill_stateReg_string = "INIT ";
      MmuPlugin_logic_refill_enumDef_CMD_0 : MmuPlugin_logic_refill_stateReg_string = "CMD_0";
      MmuPlugin_logic_refill_enumDef_CMD_1 : MmuPlugin_logic_refill_stateReg_string = "CMD_1";
      MmuPlugin_logic_refill_enumDef_RSP_0 : MmuPlugin_logic_refill_stateReg_string = "RSP_0";
      MmuPlugin_logic_refill_enumDef_RSP_1 : MmuPlugin_logic_refill_stateReg_string = "RSP_1";
      default : MmuPlugin_logic_refill_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateNext)
      MmuPlugin_logic_refill_enumDef_BOOT : MmuPlugin_logic_refill_stateNext_string = "BOOT ";
      MmuPlugin_logic_refill_enumDef_IDLE : MmuPlugin_logic_refill_stateNext_string = "IDLE ";
      MmuPlugin_logic_refill_enumDef_INIT : MmuPlugin_logic_refill_stateNext_string = "INIT ";
      MmuPlugin_logic_refill_enumDef_CMD_0 : MmuPlugin_logic_refill_stateNext_string = "CMD_0";
      MmuPlugin_logic_refill_enumDef_CMD_1 : MmuPlugin_logic_refill_stateNext_string = "CMD_1";
      MmuPlugin_logic_refill_enumDef_RSP_0 : MmuPlugin_logic_refill_stateNext_string = "RSP_0";
      MmuPlugin_logic_refill_enumDef_RSP_1 : MmuPlugin_logic_refill_stateNext_string = "RSP_1";
      default : MmuPlugin_logic_refill_stateNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "BITWISE ";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "AND_1";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "JALR";
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "JALR";
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "????";
    endcase
  end
  always @(*) begin
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_BOOT : PrivilegedPlugin_logic_fsm_stateReg_string = "BOOT      ";
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : PrivilegedPlugin_logic_fsm_stateReg_string = "IDLE      ";
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : PrivilegedPlugin_logic_fsm_stateReg_string = "SETUP     ";
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : PrivilegedPlugin_logic_fsm_stateReg_string = "EPC_WRITE ";
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : PrivilegedPlugin_logic_fsm_stateReg_string = "TVAL_WRITE";
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : PrivilegedPlugin_logic_fsm_stateReg_string = "EPC_READ  ";
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : PrivilegedPlugin_logic_fsm_stateReg_string = "TVEC_READ ";
      PrivilegedPlugin_logic_fsm_enumDef_XRET : PrivilegedPlugin_logic_fsm_stateReg_string = "XRET      ";
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : PrivilegedPlugin_logic_fsm_stateReg_string = "FLUSH_CALC";
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : PrivilegedPlugin_logic_fsm_stateReg_string = "FLUSH_JUMP";
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : PrivilegedPlugin_logic_fsm_stateReg_string = "TRAP      ";
      default : PrivilegedPlugin_logic_fsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(PrivilegedPlugin_logic_fsm_stateNext)
      PrivilegedPlugin_logic_fsm_enumDef_BOOT : PrivilegedPlugin_logic_fsm_stateNext_string = "BOOT      ";
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : PrivilegedPlugin_logic_fsm_stateNext_string = "IDLE      ";
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : PrivilegedPlugin_logic_fsm_stateNext_string = "SETUP     ";
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : PrivilegedPlugin_logic_fsm_stateNext_string = "EPC_WRITE ";
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : PrivilegedPlugin_logic_fsm_stateNext_string = "TVAL_WRITE";
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : PrivilegedPlugin_logic_fsm_stateNext_string = "EPC_READ  ";
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : PrivilegedPlugin_logic_fsm_stateNext_string = "TVEC_READ ";
      PrivilegedPlugin_logic_fsm_enumDef_XRET : PrivilegedPlugin_logic_fsm_stateNext_string = "XRET      ";
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : PrivilegedPlugin_logic_fsm_stateNext_string = "FLUSH_CALC";
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : PrivilegedPlugin_logic_fsm_stateNext_string = "FLUSH_JUMP";
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : PrivilegedPlugin_logic_fsm_stateNext_string = "TRAP      ";
      default : PrivilegedPlugin_logic_fsm_stateNext_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    if(EU0_ExecutionUnitBase_pipeline_completion_0_port_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(Lsu2Plugin_setup_specialCompletion_valid) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(Lsu2Plugin_setup_sharedCompletion_valid) begin
      _zz_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_5 = 1'b0;
    if(RobPlugin_logic_completionMem_targetWrite_valid) begin
      _zz_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_6 = 1'b0;
    if(BranchContextPlugin_free_dispatchMem_writes_0_port_valid) begin
      _zz_6 = 1'b1;
    end
  end

  always @(*) begin
    DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_1 = DecoderPredictionPlugin_logic_decodePatch_rasPushUsed;
    if(when_DecoderPredictionPlugin_l212) begin
      DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_7 = 1'b0;
    if(CsrRamPlugin_logic_writeLogic_port_valid) begin
      _zz_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_8 = 1'b0;
    if(EU0_BranchPlugin_logic_branch_finalBranch_valid) begin
      _zz_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548 = 1'b0;
    if(Lsu2Plugin_logic_flush_busy) begin
      _zz_FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548 = 1'b1;
    end
  end

  always @(*) begin
    _zz_9 = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(!when_Lsu2Plugin_l1374) begin
              _zz_9 = 1'b1;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    _zz_10 = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(!when_Lsu2Plugin_l1333) begin
              _zz_10 = 1'b1;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    _zz_11 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_11 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_12 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_12 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_13 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_13 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_14 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_14 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_15 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_15 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_16 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_16 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_17 = 1'b0;
    if(when_Lsu2Plugin_l959) begin
      _zz_17 = 1'b1;
    end
  end

  always @(*) begin
    _zz_Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842 = 1'b0;
    if(when_Lsu2Plugin_l841) begin
      _zz_Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842 = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_allocation_stores_alloc_1 = Lsu2Plugin_logic_allocation_stores_alloc;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      Lsu2Plugin_logic_allocation_stores_alloc_1 = (Lsu2Plugin_logic_allocation_stores_alloc + 4'b0001);
    end
  end

  always @(*) begin
    _zz_18 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_18 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_19 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_19 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_20 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_20 = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_allocation_loads_alloc_1 = Lsu2Plugin_logic_allocation_loads_alloc;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      Lsu2Plugin_logic_allocation_loads_alloc_1 = (Lsu2Plugin_logic_allocation_loads_alloc + 4'b0001);
    end
  end

  always @(*) begin
    _zz_21 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_21 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_22 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_22 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_23 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_23 = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_onCommit_commitComb_1 = Lsu2Plugin_logic_sq_onCommit_commitComb;
    Lsu2Plugin_logic_sq_onCommit_commitComb_1 = (Lsu2Plugin_logic_sq_onCommit_commitComb + _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1);
  end

  always @(*) begin
    _zz_24 = 1'b0;
    if(Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_valid) begin
      _zz_24 = 1'b1;
    end
  end

  always @(*) begin
    _zz_25 = 1'b0;
    if(Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_valid) begin
      _zz_25 = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_onCommit_free_1 = Lsu2Plugin_logic_lq_onCommit_free;
    Lsu2Plugin_logic_lq_onCommit_free_1 = (Lsu2Plugin_logic_lq_onCommit_free + _zz_Lsu2Plugin_logic_lq_onCommit_free_1);
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_onCommit_priority_1 = Lsu2Plugin_logic_lq_onCommit_priority;
    if(Lsu2Plugin_logic_lq_onCommit_lqCommits_0) begin
      Lsu2Plugin_logic_lq_onCommit_priority_1 = ((Lsu2Plugin_logic_lq_onCommit_priority == 7'h00) ? 7'h7f : _zz_Lsu2Plugin_logic_lq_onCommit_priority_1);
    end
  end

  always @(*) begin
    HistoryPlugin_logic_update_pushes_2_stateNext_1 = HistoryPlugin_logic_update_pushes_2_stateNext;
    if(when_HistoryPlugin_l115_1) begin
      HistoryPlugin_logic_update_pushes_2_stateNext_1 = _zz_HistoryPlugin_logic_update_pushes_2_stateNext_1[23:0];
    end
  end

  always @(*) begin
    HistoryPlugin_logic_update_pushes_0_stateNext_1 = HistoryPlugin_logic_update_pushes_0_stateNext;
    if(when_HistoryPlugin_l115) begin
      HistoryPlugin_logic_update_pushes_0_stateNext_1 = _zz_HistoryPlugin_logic_update_pushes_0_stateNext_1[23:0];
    end
  end

  always @(*) begin
    HistoryPlugin_logic_onCommit_valueNext_1 = HistoryPlugin_logic_onCommit_valueNext;
    if(when_HistoryPlugin_l90) begin
      HistoryPlugin_logic_onCommit_valueNext_1 = _zz_HistoryPlugin_logic_onCommit_valueNext_1[23:0];
    end
  end

  always @(*) begin
    CommitPlugin_logic_commit_continue_1 = CommitPlugin_logic_commit_continue;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_0_enable) begin
        if(when_CommitPlugin_l211) begin
          CommitPlugin_logic_commit_continue_1 = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    _zz_26 = 1'b0;
    if(GSharePlugin_logic_mem_write_valid) begin
      _zz_26 = 1'b1;
    end
  end

  always @(*) begin
    _zz_27 = 1'b0;
    if(BtbPlugin_logic_onLearn_port_valid) begin
      _zz_27 = 1'b1;
    end
  end

  always @(*) begin
    _zz_28 = 1'b0;
    if(DecoderPredictionPlugin_logic_ras_write_valid) begin
      _zz_28 = 1'b1;
    end
  end

  always @(*) begin
    _zz_29 = 1'b0;
    if(when_BranchContextPlugin_l97) begin
      if(FrontendPlugin_allocated_ready) begin
        _zz_29 = 1'b1;
      end
    end
  end

  always @(*) begin
    BranchContextPlugin_logic_alloc_allocNext_1 = BranchContextPlugin_logic_alloc_allocNext;
    if(when_BranchContextPlugin_l97) begin
      BranchContextPlugin_logic_alloc_allocNext_1 = (BranchContextPlugin_logic_alloc_allocNext + 3'b001);
    end
  end

  always @(*) begin
    AlignerPlugin_logic_slices_remains_1 = AlignerPlugin_logic_slices_remains;
    AlignerPlugin_logic_slices_remains_1 = (AlignerPlugin_logic_slices_remains & (~ (AlignerPlugin_logic_extractors_0_valid ? AlignerPlugin_logic_extractors_0_usage : 2'b00)));
  end

  always @(*) begin
    AlignerPlugin_logic_slices_carry_1 = AlignerPlugin_logic_slices_carry;
    AlignerPlugin_logic_slices_carry_1 = (AlignerPlugin_logic_slices_carry & (~ AlignerPlugin_logic_extractors_0_usage));
  end

  always @(*) begin
    AlignerPlugin_logic_slices_used_1 = AlignerPlugin_logic_slices_used;
    AlignerPlugin_logic_slices_used_1 = (AlignerPlugin_logic_slices_used | AlignerPlugin_logic_extractors_0_usage);
  end

  always @(*) begin
    _zz_FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552 = 1'b0;
    if(FetchCachePlugin_logic_read_ctrl_redoIt) begin
      _zz_FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552 = 1'b1;
    end
  end

  always @(*) begin
    _zz_FetchPlugin_stages_2_isFlushingRoot = 1'b0;
    if(FetchCachePlugin_logic_read_ctrl_redoIt) begin
      _zz_FetchPlugin_stages_2_isFlushingRoot = 1'b1;
    end
  end

  always @(*) begin
    _zz_30 = 1'b0;
    if(FetchCachePlugin_logic_banks_0_write_valid) begin
      _zz_30 = 1'b1;
    end
  end

  always @(*) begin
    PcPlugin_logic_jump_target_1 = PcPlugin_logic_jump_target;
    if(when_PcPlugin_l57) begin
      PcPlugin_logic_jump_target_1 = (_zz_PcPlugin_logic_jump_target_1 ? BtbPlugin_setup_btbJump_payload_pc : 32'h00000000);
    end
  end

  always @(*) begin
    MmuPlugin_setup_invalidatePort_cmd_valid = 1'b0;
    if(when_CsrAccessPlugin_l183) begin
      if(!when_MmuPlugin_l218) begin
        MmuPlugin_setup_invalidatePort_cmd_valid = 1'b1;
      end
    end
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
        if(EnvCallPlugin_logic_flushes_vmaInv) begin
          MmuPlugin_setup_invalidatePort_cmd_valid = 1'b1;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    MmuPlugin_setup_invalidatePort_rsp_valid = 1'b0;
    if(when_MmuPlugin_l545) begin
      MmuPlugin_setup_invalidatePort_rsp_valid = 1'b1;
    end
  end

  assign _zz_FetchPlugin_stages_1_MMU_IO = (_zz__zz_FetchPlugin_stages_1_MMU_IO - 32'h00000001);
  always @(*) begin
    FetchCachePlugin_setup_invalidatePort_cmd_valid = 1'b0;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
        if(EnvCallPlugin_logic_flushes_fetchInv) begin
          FetchCachePlugin_setup_invalidatePort_cmd_valid = 1'b1;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_invalidatePort_rsp_valid = 1'b0;
    if(when_FetchCachePlugin_l400) begin
      FetchCachePlugin_setup_invalidatePort_rsp_valid = 1'b1;
    end
  end

  assign AlignerPlugin_setup_singleFetch = 1'b0;
  assign FrontendPlugin_decoded_isFireing = (FrontendPlugin_decoded_valid && FrontendPlugin_decoded_ready);
  assign FrontendPlugin_allocated_isFireing = (FrontendPlugin_allocated_valid && FrontendPlugin_allocated_ready);
  always @(*) begin
    DecoderPlugin_setup_trapHalt = 1'b0;
    if(PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt) begin
      DecoderPlugin_setup_trapHalt = 1'b1;
    end
  end

  always @(*) begin
    DecoderPlugin_setup_trapRaise = 1'b0;
    if(when_PrivilegedPlugin_l679) begin
      DecoderPlugin_setup_trapRaise = 1'b1;
    end
  end

  assign DecoderPlugin_setup_debugEnter_0 = 1'b0;
  always @(*) begin
    Lsu2Plugin_setup_postCommitBusy = 1'b0;
    if(when_Lsu2Plugin_l572) begin
      Lsu2Plugin_setup_postCommitBusy = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_flushPort_cmd_valid = 1'b0;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
        Lsu2Plugin_setup_flushPort_cmd_valid = 1'b1;
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_flushPort_cmd_payload_withFree = 1'bx;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
        Lsu2Plugin_setup_flushPort_cmd_payload_withFree = EnvCallPlugin_logic_flushes_flushData;
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_flushPort_rsp_valid = 1'b0;
    if(when_Lsu2Plugin_l1553) begin
      if(when_Lsu2Plugin_l1569) begin
        Lsu2Plugin_setup_flushPort_rsp_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    PrivilegedPlugin_setup_jump_valid = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
        PrivilegedPlugin_setup_jump_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
        PrivilegedPlugin_setup_jump_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_setup_jump_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_jump_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
        PrivilegedPlugin_setup_jump_payload_pc = PrivilegedPlugin_logic_readed;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
        PrivilegedPlugin_setup_jump_payload_pc = PrivilegedPlugin_logic_readed;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_setup_jump_payload_pc = PrivilegedPlugin_logic_readed;
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_setup_withMachinePrivilege = (2'b11 <= PrivilegedPlugin_setup_privilege);
  assign PrivilegedPlugin_setup_withSupervisorPrivilege = (2'b01 <= PrivilegedPlugin_setup_privilege);
  always @(*) begin
    PrivilegedPlugin_setup_xretAwayFromMachine = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
        if(when_PrivilegedPlugin_l959) begin
          PrivilegedPlugin_setup_xretAwayFromMachine = 1'b1;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_trapEvent = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_setup_trapEvent = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_redoTriggered = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
        if(!when_PrivilegedPlugin_l773) begin
          case(PrivilegedPlugin_logic_reschedule_payload_cause)
            4'b1001 : begin
            end
            4'b1010 : begin
              PrivilegedPlugin_setup_redoTriggered = 1'b1;
            end
            4'b1000 : begin
            end
            default : begin
            end
          endcase
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_setup_setFpDirty = 1'b0;
  assign PrivilegedPlugin_setup_isFpuEnabled = 1'b0;
  always @(*) begin
    EU0_CsrAccessPlugin_setup_onDecodeTrap = 1'b0;
    if(when_PrivilegedPlugin_l165) begin
      EU0_CsrAccessPlugin_setup_onDecodeTrap = 1'b1;
    end
    if(when_CsrAccessPlugin_l183) begin
      if(when_MmuPlugin_l218) begin
        EU0_CsrAccessPlugin_setup_onDecodeTrap = 1'b1;
      end
    end
  end

  always @(*) begin
    EU0_CsrAccessPlugin_setup_onDecodeFlushPipeline = 1'b0;
    if(when_CsrAccessPlugin_l183) begin
      if(!when_MmuPlugin_l218) begin
        EU0_CsrAccessPlugin_setup_onDecodeFlushPipeline = 1'b1;
      end
    end
  end

  always @(*) begin
    EU0_CsrAccessPlugin_setup_onReadHalt = 1'b0;
    if(when_CsrAccessPlugin_l272) begin
      EU0_CsrAccessPlugin_setup_onReadHalt = 1'b1;
    end
  end

  always @(*) begin
    EU0_CsrAccessPlugin_setup_onWriteHalt = 1'b0;
    if(when_CsrAccessPlugin_l342) begin
      EU0_CsrAccessPlugin_setup_onWriteHalt = 1'b1;
    end
  end

  assign EU0_CsrAccessPlugin_setup_onWriteFlushPipeline = 1'b0;
  assign clint_awready = clintCtrl_io_bus_aw_ready;
  assign clint_wready = clintCtrl_io_bus_w_ready;
  assign clint_bvalid = clintCtrl_io_bus_b_valid;
  assign clint_bresp = clintCtrl_io_bus_b_payload_resp;
  assign clint_arready = clintCtrl_io_bus_ar_ready;
  assign clint_rvalid = clintCtrl_io_bus_r_valid;
  assign clint_rdata = clintCtrl_io_bus_r_payload_data;
  assign clint_rresp = clintCtrl_io_bus_r_payload_resp;
  assign plic_awready = plicCtrl_io_bus_aw_ready;
  assign plic_wready = plicCtrl_io_bus_w_ready;
  assign plic_bvalid = plicCtrl_io_bus_b_valid;
  assign plic_bresp = plicCtrl_io_bus_b_payload_resp;
  assign plic_arready = plicCtrl_io_bus_ar_ready;
  assign plic_rvalid = plicCtrl_io_bus_r_valid;
  assign plic_rdata = plicCtrl_io_bus_r_payload_data;
  assign plic_rresp = plicCtrl_io_bus_r_payload_resp;
  assign plicCtrl_io_sources = (plicInterrupts >>> 1'd1);
  assign iBusAxi_arvalid = FetchCachePlugin_mem_cmd_valid;
  assign iBusAxi_araddr = FetchCachePlugin_mem_cmd_payload_address;
  assign iBusAxi_arprot = 3'b110;
  assign iBusAxi_arlen = 8'h0f;
  assign iBusAxi_arsize = 3'b010;
  assign iBusAxi_arburst = 2'b01;
  assign FetchCachePlugin_mem_cmd_ready = iBusAxi_arready;
  assign FetchCachePlugin_mem_rsp_valid = iBusAxi_rvalid;
  assign FetchCachePlugin_mem_rsp_payload_data = iBusAxi_rdata;
  assign FetchCachePlugin_mem_rsp_payload_error = (! (iBusAxi_rresp == 2'b00));
  assign iBusAxi_rready = 1'b1;
  assign FetchPlugin_stages_1_isFireing = (FetchPlugin_stages_1_valid && FetchPlugin_stages_1_ready);
  assign when_Stage_l170 = (FetchPlugin_stages_1_ready || FetchPlugin_stages_1_isFlushed);
  assign FetchPlugin_stages_1_isFirstCycle = (FetchPlugin_stages_1_valid && (! _zz_FetchPlugin_stages_1_isFirstCycle));
  assign _zz_PcPlugin_logic_jump_oh = {BtbPlugin_setup_btbJump_valid,{FetchCachePlugin_setup_redoJump_valid,{AlignerPlugin_setup_sequenceJump_valid,{DecoderPredictionPlugin_setup_decodeJump_valid,{CommitPlugin_setup_jump_valid,PrivilegedPlugin_setup_jump_valid}}}}};
  assign _zz_PcPlugin_logic_jump_oh_1 = _zz_PcPlugin_logic_jump_oh[0];
  assign _zz_PcPlugin_logic_jump_oh_2 = _zz_PcPlugin_logic_jump_oh[1];
  assign _zz_PcPlugin_logic_jump_oh_3 = _zz_PcPlugin_logic_jump_oh[2];
  assign _zz_PcPlugin_logic_jump_oh_4 = _zz_PcPlugin_logic_jump_oh[3];
  assign _zz_PcPlugin_logic_jump_oh_5 = _zz_PcPlugin_logic_jump_oh[4];
  always @(*) begin
    _zz_PcPlugin_logic_jump_oh_6[0] = (_zz_PcPlugin_logic_jump_oh_1 && (! 1'b0));
    _zz_PcPlugin_logic_jump_oh_6[1] = (_zz_PcPlugin_logic_jump_oh_2 && (! _zz_PcPlugin_logic_jump_oh_1));
    _zz_PcPlugin_logic_jump_oh_6[2] = (_zz_PcPlugin_logic_jump_oh_3 && (! (|{_zz_PcPlugin_logic_jump_oh_2,_zz_PcPlugin_logic_jump_oh_1})));
    _zz_PcPlugin_logic_jump_oh_6[3] = (_zz_PcPlugin_logic_jump_oh_4 && (! (|{_zz_PcPlugin_logic_jump_oh_3,{_zz_PcPlugin_logic_jump_oh_2,_zz_PcPlugin_logic_jump_oh_1}})));
    _zz_PcPlugin_logic_jump_oh_6[4] = (_zz_PcPlugin_logic_jump_oh_5 && (! _zz_PcPlugin_logic_jump_oh_7));
    _zz_PcPlugin_logic_jump_oh_6[5] = (_zz_PcPlugin_logic_jump_oh[5] && (! (_zz_PcPlugin_logic_jump_oh_5 || _zz_PcPlugin_logic_jump_oh_7)));
  end

  assign _zz_PcPlugin_logic_jump_oh_7 = (|{_zz_PcPlugin_logic_jump_oh_4,{_zz_PcPlugin_logic_jump_oh_3,{_zz_PcPlugin_logic_jump_oh_2,_zz_PcPlugin_logic_jump_oh_1}}});
  assign PcPlugin_logic_jump_oh = _zz_PcPlugin_logic_jump_oh_6;
  assign PcPlugin_logic_jump_target = ((((PcPlugin_logic_jump_oh[0] ? PrivilegedPlugin_setup_jump_payload_pc : 32'h00000000) | (PcPlugin_logic_jump_oh[1] ? CommitPlugin_setup_jump_payload_pc : 32'h00000000)) | ((PcPlugin_logic_jump_oh[2] ? DecoderPredictionPlugin_setup_decodeJump_payload_pc : 32'h00000000) | (PcPlugin_logic_jump_oh[3] ? AlignerPlugin_setup_sequenceJump_payload_pc : 32'h00000000))) | (PcPlugin_logic_jump_oh[4] ? FetchCachePlugin_setup_redoJump_payload_pc : 32'h00000000));
  assign _zz_PcPlugin_logic_jump_target_1 = PcPlugin_logic_jump_oh[5];
  assign when_PcPlugin_l57 = (|_zz_PcPlugin_logic_jump_target_1);
  assign PcPlugin_logic_jump_pcLoad_valid = (|{PrivilegedPlugin_setup_jump_valid,{CommitPlugin_setup_jump_valid,{BtbPlugin_setup_btbJump_valid,{DecoderPredictionPlugin_setup_decodeJump_valid,{AlignerPlugin_setup_sequenceJump_valid,FetchCachePlugin_setup_redoJump_valid}}}}});
  assign PcPlugin_logic_jump_pcLoad_payload_pc = PcPlugin_logic_jump_target_1;
  assign FetchCachePlugin_logic_banks_0_read_rsp = FetchCachePlugin_logic_banks_0_mem_spinal_port1;
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_0 = FetchCachePlugin_logic_banks_0_read_rsp;
  always @(*) begin
    FetchCachePlugin_logic_waysWrite_mask = 1'b0;
    if(when_FetchCachePlugin_l383) begin
      FetchCachePlugin_logic_waysWrite_mask = 1'b1;
    end
    if(FetchCachePlugin_logic_invalidate_done) begin
      if(FetchCachePlugin_logic_refill_fire) begin
        FetchCachePlugin_logic_waysWrite_mask[0] = 1'b1;
      end
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_waysWrite_address = 2'bxx;
    if(when_FetchCachePlugin_l383) begin
      FetchCachePlugin_logic_waysWrite_address = FetchCachePlugin_logic_invalidate_counter[1:0];
    end
    if(FetchCachePlugin_logic_invalidate_done) begin
      FetchCachePlugin_logic_waysWrite_address = FetchCachePlugin_logic_refill_address[7 : 6];
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_waysWrite_tag_loaded = 1'bx;
    if(when_FetchCachePlugin_l383) begin
      FetchCachePlugin_logic_waysWrite_tag_loaded = 1'b0;
    end
    if(FetchCachePlugin_logic_invalidate_done) begin
      FetchCachePlugin_logic_waysWrite_tag_loaded = 1'b1;
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_waysWrite_tag_error = 1'bx;
    if(FetchCachePlugin_logic_invalidate_done) begin
      FetchCachePlugin_logic_waysWrite_tag_error = (FetchCachePlugin_logic_refill_hadError || FetchCachePlugin_mem_rsp_payload_error);
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_waysWrite_tag_address = 24'bxxxxxxxxxxxxxxxxxxxxxxxx;
    if(FetchCachePlugin_logic_invalidate_done) begin
      FetchCachePlugin_logic_waysWrite_tag_address = FetchCachePlugin_logic_refill_address[31 : 8];
    end
  end

  assign _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded = FetchCachePlugin_logic_ways_0_mem_spinal_port1;
  assign FetchCachePlugin_logic_ways_0_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded[0];
  assign FetchCachePlugin_logic_ways_0_read_rsp_error = _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded[1];
  assign FetchCachePlugin_logic_ways_0_read_rsp_address = _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded[25 : 2];
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_loaded = FetchCachePlugin_logic_ways_0_read_rsp_loaded;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_error = FetchCachePlugin_logic_ways_0_read_rsp_error;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_address = FetchCachePlugin_logic_ways_0_read_rsp_address;
  always @(*) begin
    FetchCachePlugin_logic_invalidate_canStart = 1'b1;
    if(when_FetchCachePlugin_l396) begin
      FetchCachePlugin_logic_invalidate_canStart = 1'b0;
    end
    if(FetchCachePlugin_logic_refill_valid) begin
      FetchCachePlugin_logic_invalidate_canStart = 1'b0;
    end
  end

  assign FetchCachePlugin_logic_invalidate_done = FetchCachePlugin_logic_invalidate_counter[2];
  assign when_FetchCachePlugin_l379 = (! FetchCachePlugin_logic_invalidate_done);
  assign when_FetchCachePlugin_l383 = (! FetchCachePlugin_logic_invalidate_done);
  assign FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l389 = ((! FetchCachePlugin_logic_invalidate_done) || FetchCachePlugin_logic_invalidate_requested);
  assign when_FetchCachePlugin_l391 = (FetchCachePlugin_logic_invalidate_requested && FetchCachePlugin_logic_invalidate_canStart);
  assign when_FetchCachePlugin_l396 = (|{FetchPlugin_stages_2_valid,FetchPlugin_stages_1_valid});
  assign when_FetchCachePlugin_l400 = (FetchCachePlugin_logic_invalidate_done && (! FetchCachePlugin_logic_invalidate_done_regNext));
  always @(*) begin
    FetchCachePlugin_logic_refill_start_valid = 1'b0;
    if(FetchPlugin_stages_2_valid) begin
      if(!FetchPlugin_stages_2_MMU_REDO) begin
        if(when_FetchCachePlugin_l562) begin
          FetchCachePlugin_logic_refill_start_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_refill_fire = 1'b0;
    if(FetchCachePlugin_mem_rsp_valid) begin
      if(when_FetchCachePlugin_l470) begin
        FetchCachePlugin_logic_refill_fire = 1'b1;
      end
    end
  end

  assign when_FetchCachePlugin_l422 = (! FetchCachePlugin_logic_refill_valid);
  assign FetchCachePlugin_mem_cmd_fire = (FetchCachePlugin_mem_cmd_valid && FetchCachePlugin_mem_cmd_ready);
  assign FetchCachePlugin_mem_cmd_valid = (FetchCachePlugin_logic_refill_valid && (! FetchCachePlugin_logic_refill_cmdSent));
  assign FetchCachePlugin_mem_cmd_payload_address = {FetchCachePlugin_logic_refill_address[31 : 6],6'h00};
  assign FetchCachePlugin_mem_cmd_payload_io = FetchCachePlugin_logic_refill_isIo;
  assign when_Utils_l578 = (! FetchCachePlugin_logic_refill_valid);
  always @(*) begin
    FetchCachePlugin_logic_refill_randomWay_willIncrement = 1'b0;
    if(when_Utils_l578) begin
      FetchCachePlugin_logic_refill_randomWay_willIncrement = 1'b1;
    end
  end

  assign FetchCachePlugin_logic_refill_randomWay_willClear = 1'b0;
  assign FetchCachePlugin_logic_refill_randomWay_willOverflowIfInc = 1'b1;
  assign FetchCachePlugin_logic_refill_randomWay_willOverflow = (FetchCachePlugin_logic_refill_randomWay_willOverflowIfInc && FetchCachePlugin_logic_refill_randomWay_willIncrement);
  assign FetchCachePlugin_logic_banks_0_write_valid = (FetchCachePlugin_mem_rsp_valid && 1'b1);
  assign FetchCachePlugin_logic_banks_0_write_payload_address = {FetchCachePlugin_logic_refill_address[7 : 6],FetchCachePlugin_logic_refill_wordIndex};
  assign FetchCachePlugin_logic_banks_0_write_payload_data = FetchCachePlugin_mem_rsp_payload_data;
  assign FetchCachePlugin_mem_rsp_ready = 1'b1;
  assign when_FetchCachePlugin_l470 = (FetchCachePlugin_logic_refill_wordIndex == 4'b1111);
  assign FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l476 = FetchCachePlugin_logic_refill_valid;
  assign FetchCachePlugin_logic_banks_0_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_banks_0_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[7 : 2];
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_0 = FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_0[31 : 0];
  assign FetchPlugin_stages_2_Fetch_WORD = (FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_0 ? FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_0 : 32'h00000000);
  assign FetchCachePlugin_logic_ways_0_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_ways_0_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[7 : 6];
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_0 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0[31 : 8]) && FetchPlugin_stages_1_MMU_WAYS_OH[0]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_1 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1[31 : 8]) && FetchPlugin_stages_1_MMU_WAYS_OH[1]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_2 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2[31 : 8]) && FetchPlugin_stages_1_MMU_WAYS_OH[2]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_3 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3[31 : 8]) && FetchPlugin_stages_1_MMU_WAYS_OH[3]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_4 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4[31 : 8]) && FetchPlugin_stages_1_MMU_WAYS_OH[4]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_5 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5[31 : 8]) && FetchPlugin_stages_1_MMU_WAYS_OH[5]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_translatedHits = (|{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_5,{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_4,{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_3,{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_2,{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_1,FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_0}}}}});
  assign FetchCachePlugin_logic_read_onWays_0_hits_bypassHits = (FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == _zz_FetchCachePlugin_logic_read_onWays_0_hits_bypassHits);
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_0 = ((FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION ? FetchCachePlugin_logic_read_onWays_0_hits_bypassHits : FetchCachePlugin_logic_read_onWays_0_hits_translatedHits) && FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_loaded);
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HIT = (|FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_0);
  always @(*) begin
    FetchCachePlugin_logic_plru_write_valid = 1'b0;
    if(!FetchCachePlugin_logic_read_ctrl_redoIt) begin
      if(FetchPlugin_stages_2_isFireing) begin
        FetchCachePlugin_logic_plru_write_valid = 1'b1;
      end
    end
    if(when_FetchCachePlugin_l593) begin
      FetchCachePlugin_logic_plru_write_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_plru_write_payload_address = FetchPlugin_stages_2_Fetch_FETCH_PC[7 : 6];
    if(when_FetchCachePlugin_l593) begin
      FetchCachePlugin_logic_plru_write_payload_address = FetchCachePlugin_logic_invalidate_counter[1:0];
    end
  end

  always @(*) begin
    FetchCachePlugin_setup_redoJump_valid = 1'b0;
    if(FetchCachePlugin_logic_read_ctrl_redoIt) begin
      FetchCachePlugin_setup_redoJump_valid = 1'b1;
    end
  end

  assign FetchCachePlugin_setup_redoJump_payload_pc = FetchPlugin_stages_2_Fetch_FETCH_PC;
  assign FetchPlugin_stages_2_Fetch_WORD_FAULT = (((|(FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_0 & FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_error)) || FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE) || FetchPlugin_stages_2_MMU_ACCESS_FAULT);
  assign FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE = (FetchPlugin_stages_2_MMU_PAGE_FAULT || (! FetchPlugin_stages_2_MMU_ALLOW_EXECUTE));
  always @(*) begin
    FetchCachePlugin_logic_read_ctrl_redoIt = 1'b0;
    if(FetchPlugin_stages_2_valid) begin
      if(FetchPlugin_stages_2_MMU_REDO) begin
        FetchCachePlugin_logic_read_ctrl_redoIt = 1'b1;
      end else begin
        if(when_FetchCachePlugin_l562) begin
          FetchCachePlugin_logic_read_ctrl_redoIt = 1'b1;
        end
      end
    end
  end

  assign FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552 = _zz_FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552;
  assign FetchPlugin_stages_2_isFireing = (FetchPlugin_stages_2_valid && FetchPlugin_stages_2_ready);
  assign when_FetchCachePlugin_l562 = (((! FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE) && (! FetchPlugin_stages_2_MMU_ACCESS_FAULT)) && (! FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HIT));
  assign FetchCachePlugin_logic_refill_start_address = FetchPlugin_stages_2_MMU_TRANSLATED;
  assign FetchCachePlugin_logic_refill_start_isIo = FetchPlugin_stages_2_MMU_IO;
  assign FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l583 = (! FetchCachePlugin_logic_translationPort_wake);
  assign FetchCachePlugin_setup_historyJump_valid = FetchCachePlugin_setup_redoJump_valid;
  assign FetchCachePlugin_setup_historyJump_payload_history = FetchPlugin_stages_2_BRANCH_HISTORY;
  assign when_FetchCachePlugin_l593 = ((! FetchCachePlugin_logic_invalidate_done) && FetchCachePlugin_logic_invalidate_firstEver);
  assign AlignerPlugin_logic_ignoreInput = AlignerPlugin_setup_s2m_isFlushingRoot;
  assign AlignerPlugin_logic_isInputValid = (AlignerPlugin_setup_s2m_valid && (! AlignerPlugin_logic_ignoreInput));
  assign FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT = 1'b1;
  always @(*) begin
    AlignerPlugin_setup_s2m_MASK_BACK = 1'b1;
    if(when_AlignerPlugin_l98) begin
      AlignerPlugin_setup_s2m_MASK_BACK = 1'b1;
    end
  end

  assign when_AlignerPlugin_l98 = (! AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID);
  assign _zz_AlignerPlugin_logic_slices_data_0 = {AlignerPlugin_setup_s2m_Fetch_WORD,AlignerPlugin_logic_buffer_data};
  assign AlignerPlugin_logic_slices_data_0 = _zz_AlignerPlugin_logic_slices_data_0[31 : 0];
  assign AlignerPlugin_logic_slices_data_1 = _zz_AlignerPlugin_logic_slices_data_0[63 : 32];
  assign AlignerPlugin_logic_slices_carry = {(AlignerPlugin_logic_isInputValid ? AlignerPlugin_setup_s2m_MASK_FRONT : 1'b0),AlignerPlugin_logic_buffer_mask};
  assign AlignerPlugin_logic_slices_remains = AlignerPlugin_logic_slices_carry;
  assign AlignerPlugin_logic_slices_used = 2'b00;
  assign AlignerPlugin_logic_decoders_0_usage = 2'b01;
  assign AlignerPlugin_logic_decoders_0_notEnoughData = 1'b0;
  assign AlignerPlugin_logic_decoders_0_pastPrediction = 1'b0;
  assign AlignerPlugin_logic_decoders_0_usable = ((! AlignerPlugin_logic_decoders_0_notEnoughData) && (! AlignerPlugin_logic_decoders_0_pastPrediction));
  assign AlignerPlugin_logic_decoders_1_usage = 2'b10;
  assign AlignerPlugin_logic_decoders_1_notEnoughData = 1'b0;
  assign AlignerPlugin_logic_decoders_1_pastPrediction = 1'b0;
  assign AlignerPlugin_logic_decoders_1_usable = ((! AlignerPlugin_logic_decoders_1_notEnoughData) && (! AlignerPlugin_logic_decoders_1_pastPrediction));
  assign _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_maskOh = AlignerPlugin_logic_slices_carry[1 : 0];
  assign _zz_AlignerPlugin_logic_extractors_0_maskOh_1 = _zz_AlignerPlugin_logic_extractors_0_maskOh[0];
  always @(*) begin
    _zz_AlignerPlugin_logic_extractors_0_maskOh_2[0] = (_zz_AlignerPlugin_logic_extractors_0_maskOh_1 && (! 1'b0));
    _zz_AlignerPlugin_logic_extractors_0_maskOh_2[1] = (_zz_AlignerPlugin_logic_extractors_0_maskOh[1] && (! _zz_AlignerPlugin_logic_extractors_0_maskOh_1));
  end

  assign AlignerPlugin_logic_extractors_0_maskOh = _zz_AlignerPlugin_logic_extractors_0_maskOh_2;
  assign _zz_AlignerPlugin_logic_extractors_0_usage = AlignerPlugin_logic_extractors_0_maskOh[0];
  assign _zz_AlignerPlugin_logic_extractors_0_usage_1 = AlignerPlugin_logic_extractors_0_maskOh[1];
  assign AlignerPlugin_logic_extractors_0_usage = ((_zz_AlignerPlugin_logic_extractors_0_usage ? AlignerPlugin_logic_decoders_0_usage : 2'b00) | (_zz_AlignerPlugin_logic_extractors_0_usage_1 ? AlignerPlugin_logic_decoders_1_usage : 2'b00));
  assign AlignerPlugin_logic_extractors_0_usable = _zz_AlignerPlugin_logic_extractors_0_usable[0];
  assign AlignerPlugin_logic_extractors_0_slice0 = ((_zz_AlignerPlugin_logic_extractors_0_usage ? AlignerPlugin_logic_slices_data_0 : 32'h00000000) | (_zz_AlignerPlugin_logic_extractors_0_usage_1 ? AlignerPlugin_logic_slices_data_1 : 32'h00000000));
  assign AlignerPlugin_logic_extractors_0_valid = ((|AlignerPlugin_logic_slices_carry[1 : 0]) && AlignerPlugin_logic_extractors_0_usable);
  assign FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_0 = AlignerPlugin_logic_extractors_0_slice0;
  assign FrontendPlugin_aligned_Frontend_MASK_ALIGNED_0 = AlignerPlugin_logic_extractors_0_valid;
  assign AlignerPlugin_logic_extractors_0_bufferPredictionLast = 1'b1;
  assign AlignerPlugin_logic_extractors_0_inputPredictionLast = 1'b1;
  assign AlignerPlugin_logic_extractors_0_lastWord = (|AlignerPlugin_logic_extractors_0_maskOh[1 : 1]);
  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0 = ((AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID && (! _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0)) && AlignerPlugin_logic_extractors_0_inputPredictionLast);
    end else begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0 = (AlignerPlugin_logic_buffer_branchValid && AlignerPlugin_logic_extractors_0_bufferPredictionLast);
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_0 = AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT;
    end else begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_0 = AlignerPlugin_logic_buffer_branchPcNext;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_BRANCH_HISTORY_0 = AlignerPlugin_setup_s2m_BRANCH_HISTORY;
    end else begin
      FrontendPlugin_aligned_BRANCH_HISTORY_0 = AlignerPlugin_logic_buffer_wordContexts_0;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_0 = AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID;
    end else begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_0 = AlignerPlugin_logic_buffer_wordContexts_1;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_0 = AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE;
    end else begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_0 = AlignerPlugin_logic_buffer_wordContexts_3;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_GSHARE_COUNTER_0_0 = AlignerPlugin_setup_s2m_GSHARE_COUNTER_0;
    end else begin
      FrontendPlugin_aligned_GSHARE_COUNTER_0_0 = AlignerPlugin_logic_buffer_wordContexts_4_0;
    end
  end

  assign _zz_AlignerPlugin_logic_extractors_0_sliceOffset = AlignerPlugin_logic_extractors_0_maskOh[1];
  assign AlignerPlugin_logic_extractors_0_sliceOffset = _zz_AlignerPlugin_logic_extractors_0_sliceOffset;
  assign AlignerPlugin_logic_extractors_0_firstWord = AlignerPlugin_logic_extractors_0_sliceOffset[0];
  assign AlignerPlugin_logic_extractors_0_pcWord = _zz_AlignerPlugin_logic_extractors_0_pcWord;
  assign FrontendPlugin_aligned_PC_0 = {_zz_FrontendPlugin_aligned_PC_0,2'b00};
  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_firstWord) begin
      FrontendPlugin_aligned_FETCH_ID_0 = AlignerPlugin_setup_s2m_FETCH_ID;
    end else begin
      FrontendPlugin_aligned_FETCH_ID_0 = AlignerPlugin_logic_buffer_firstWordContexts_0;
    end
  end

  always @(*) begin
    FrontendPlugin_aligned_Frontend_FETCH_FAULT_0 = 1'b0;
    if(when_AlignerPlugin_l230) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_0 = 1'b1;
    end
    if(when_AlignerPlugin_l235) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_0 = 1'b1;
    end
  end

  always @(*) begin
    FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0 = 1'bx;
    if(when_AlignerPlugin_l230) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0 = AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE;
    end
    if(when_AlignerPlugin_l235) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0 = AlignerPlugin_logic_buffer_fault_page;
    end
  end

  assign when_AlignerPlugin_l230 = ((AlignerPlugin_logic_extractors_0_firstWord || AlignerPlugin_logic_extractors_0_lastWord) && AlignerPlugin_setup_s2m_Fetch_WORD_FAULT);
  assign when_AlignerPlugin_l235 = (((! AlignerPlugin_logic_extractors_0_firstWord) || (! AlignerPlugin_logic_extractors_0_lastWord)) && AlignerPlugin_logic_buffer_fault);
  assign FrontendPlugin_aligned_isFireing = (FrontendPlugin_aligned_valid && FrontendPlugin_aligned_ready);
  assign AlignerPlugin_logic_fireOutput = FrontendPlugin_aligned_isFireing;
  assign AlignerPlugin_logic_fireInput = ((AlignerPlugin_logic_isInputValid && (AlignerPlugin_logic_buffer_mask == 1'b0)) || (AlignerPlugin_logic_fireOutput && (AlignerPlugin_logic_slices_remains_1[0 : 0] == 1'b0)));
  assign AlignerPlugin_logic_postMask = (_zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0 ? 1'b1 : AlignerPlugin_setup_s2m_MASK_BACK);
  assign when_AlignerPlugin_l264 = (AlignerPlugin_setup_s2m_ready || AlignerPlugin_setup_s2m_isFlushed);
  assign _zz_FetchPlugin_stages_1_isFlushingRoot = (_zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0 && (! AlignerPlugin_logic_correctionSent));
  assign AlignerPlugin_setup_sequenceJump_valid = (_zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0 && (! AlignerPlugin_logic_correctionSent));
  assign AlignerPlugin_setup_sequenceJump_payload_pc = AlignerPlugin_setup_s2m_Fetch_FETCH_PC_INC;
  assign FrontendPlugin_aligned_valid = AlignerPlugin_logic_extractors_0_valid;
  assign AlignerPlugin_setup_s2m_haltRequest_AlignerPlugin_l270 = (! AlignerPlugin_logic_fireInput);
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_0 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_0;
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_0 = 1'b0;
  assign integer_RfAllocationPlugin_logic_pop_blocked = (! integer_RfAllocationPlugin_logic_allocator_io_pop_ready);
  assign FrontendPlugin_allocated_haltRequest_RfAllocationPlugin_l55 = integer_RfAllocationPlugin_logic_pop_blocked;
  assign when_RfAllocationPlugin_l63 = 1'b1;
  assign integer_RfAllocationPlugin_logic_allocator_io_pop_mask[0] = ((FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0 && FrontendPlugin_allocated_WRITE_RD_0) && when_RfAllocationPlugin_l63);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RD_0 = 6'bxxxxxx;
    if(when_RfAllocationPlugin_l63) begin
      FrontendPlugin_allocated_PHYS_RD_0 = integer_RfAllocationPlugin_logic_allocator_io_pop_values_0;
    end
  end

  assign BranchContextPlugin_logic_ptr_occupancy = (BranchContextPlugin_logic_ptr_alloc - BranchContextPlugin_logic_ptr_free);
  assign BranchContextPlugin_logic_alloc_allocNext = BranchContextPlugin_logic_ptr_alloc;
  always @(*) begin
    BranchContextPlugin_logic_alloc_full = 1'b0;
    if(when_BranchContextPlugin_l110) begin
      BranchContextPlugin_logic_alloc_full = 1'b1;
    end
  end

  assign FrontendPlugin_allocated_BRANCH_ID_0 = BranchContextPlugin_logic_alloc_allocNext[1:0];
  assign when_BranchContextPlugin_l97 = ((FrontendPlugin_allocated_valid && FrontendPlugin_allocated_BRANCH_SEL_0) && FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0);
  assign when_BranchContextPlugin_l110 = (3'b011 < BranchContextPlugin_logic_ptr_occupancy);
  assign FrontendPlugin_allocated_haltRequest_BranchContextPlugin_l111 = BranchContextPlugin_logic_alloc_full;
  always @(*) begin
    DecoderPredictionPlugin_logic_ras_ptr_pushIt = 1'b0;
    if(when_DecoderPredictionPlugin_l212) begin
      DecoderPredictionPlugin_logic_ras_ptr_pushIt = 1'b1;
    end
    if(when_DecoderPredictionPlugin_l243) begin
      DecoderPredictionPlugin_logic_ras_ptr_pushIt = 1'b0;
    end
  end

  always @(*) begin
    DecoderPredictionPlugin_logic_ras_ptr_popIt = 1'b0;
    if(when_DecoderPredictionPlugin_l219) begin
      DecoderPredictionPlugin_logic_ras_ptr_popIt = 1'b1;
    end
    if(when_DecoderPredictionPlugin_l244) begin
      DecoderPredictionPlugin_logic_ras_ptr_popIt = 1'b0;
    end
  end

  assign DecoderPredictionPlugin_logic_ras_read = DecoderPredictionPlugin_logic_ras_mem_stack_spinal_port0;
  assign DecoderPredictionPlugin_logic_ras_write_valid = DecoderPredictionPlugin_logic_ras_ptr_pushIt;
  assign DecoderPredictionPlugin_logic_ras_write_payload_address = DecoderPredictionPlugin_logic_ras_ptr_push;
  always @(*) begin
    DecoderPredictionPlugin_logic_ras_write_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_DecoderPredictionPlugin_l212) begin
      if(when_DecoderPredictionPlugin_l213) begin
        DecoderPredictionPlugin_logic_ras_write_payload_data = FrontendPlugin_serialized_PC_INC_0;
      end
    end
  end

  assign BtbPlugin_logic_onLearn_hash = BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[17 : 2];
  assign BtbPlugin_logic_onLearn_port_valid = BranchContextPlugin_setup_learnValid;
  assign BtbPlugin_logic_onLearn_port_payload_address = _zz_BtbPlugin_logic_onLearn_port_payload_address[2:0];
  assign BtbPlugin_logic_onLearn_port_payload_data_hash = BtbPlugin_logic_onLearn_hash;
  assign BtbPlugin_logic_onLearn_port_payload_data_pcTarget = BranchContextPlugin_learn_BRANCH_FINAL_pcTarget;
  assign BtbPlugin_logic_onLearn_port_payload_data_isBranch = BranchContextPlugin_free_learn_Prediction_IS_BRANCH;
  assign BtbPlugin_logic_readCmd_entryAddress = _zz_BtbPlugin_logic_readCmd_entryAddress[2:0];
  assign _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash = BtbPlugin_logic_mem_spinal_port1;
  assign FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash = _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash[15 : 0];
  assign FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_pcTarget = _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash[47 : 16];
  assign FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_isBranch = _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash[48];
  assign BtbPlugin_logic_hitCalc_postPcPrediction = 1'b0;
  assign FetchPlugin_stages_1_BtbPlugin_logic_HIT = ((FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash == FetchPlugin_stages_1_Fetch_FETCH_PC[17 : 2]) && (! BtbPlugin_logic_hitCalc_postPcPrediction));
  assign BtbPlugin_logic_applyIt_prediction = FetchPlugin_stages_1_GSHARE_COUNTER_0[1];
  assign BtbPlugin_logic_applyIt_needIt = ((FetchPlugin_stages_1_valid && FetchPlugin_stages_1_BtbPlugin_logic_HIT) && (! (FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_isBranch && (! BtbPlugin_logic_applyIt_prediction))));
  assign when_BtbPlugin_l109 = (FetchPlugin_stages_1_ready || FetchPlugin_stages_1_isFlushed);
  assign BtbPlugin_logic_applyIt_doIt = (BtbPlugin_logic_applyIt_needIt && (! BtbPlugin_logic_applyIt_correctionSent));
  assign BtbPlugin_setup_btbJump_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_setup_btbJump_payload_pc = FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_pcTarget;
  assign FetchPlugin_stages_1_Prediction_WORD_BRANCH_VALID = BtbPlugin_logic_applyIt_needIt;
  assign FetchPlugin_stages_1_Prediction_WORD_BRANCH_PC_NEXT = FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_pcTarget;
  assign BtbPlugin_setup_historyPush_flush = (((FetchPlugin_stages_1_valid && FetchPlugin_stages_1_BtbPlugin_logic_HIT) && FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_isBranch) && (! BtbPlugin_logic_applyIt_correctionSent));
  assign BtbPlugin_setup_historyPush_mask[0] = BtbPlugin_setup_historyPush_flush;
  assign BtbPlugin_setup_historyPush_taken[0] = BtbPlugin_logic_applyIt_prediction;
  assign FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALID = BtbPlugin_setup_historyPush_flush;
  assign FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALUE = BtbPlugin_logic_applyIt_prediction;
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH = FetchPlugin_stages_0_Fetch_FETCH_PC[8 : 2];
  assign FetchPlugin_stages_0_GSharePlugin_logic_HASH = ({_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[0],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[1],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[2],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[3],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[4],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[5],_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[6]}}}}}} ^ _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_1);
  assign FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_valid = GSharePlugin_logic_mem_write_valid;
  assign FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_address = GSharePlugin_logic_mem_write_payload_address;
  assign FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_0 = GSharePlugin_logic_mem_write_payload_data_0;
  always @(*) begin
    FetchPlugin_stages_1_GSHARE_COUNTER_0 = GSharePlugin_logic_mem_counter_spinal_port1[1 : 0];
    if(when_GSharePlugin_l98) begin
      FetchPlugin_stages_1_GSHARE_COUNTER_0 = FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_0;
    end
  end

  assign when_GSharePlugin_l98 = (FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_valid && (FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_address == FetchPlugin_stages_1_GSharePlugin_logic_HASH));
  assign FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_0 = FrontendPlugin_decompressed_GSHARE_COUNTER_0_0[1];
  assign _zz_GSharePlugin_logic_onLearn_hash = BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[8 : 2];
  assign GSharePlugin_logic_onLearn_hash = ({_zz_GSharePlugin_logic_onLearn_hash[0],{_zz_GSharePlugin_logic_onLearn_hash[1],{_zz_GSharePlugin_logic_onLearn_hash[2],{_zz_GSharePlugin_logic_onLearn_hash[3],{_zz_GSharePlugin_logic_onLearn_hash[4],{_zz_GSharePlugin_logic_onLearn_hash[5],_zz_GSharePlugin_logic_onLearn_hash[6]}}}}}} ^ _zz_GSharePlugin_logic_onLearn_hash_1);
  assign GSharePlugin_logic_onLearn_incrValue = (BranchContextPlugin_learn_BRANCH_FINAL_taken ? 2'b01 : 2'b11);
  always @(*) begin
    GSharePlugin_logic_onLearn_overflow = 1'b0;
    if(when_GSharePlugin_l123) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
  end

  assign GSharePlugin_logic_onLearn_updated_0 = (BranchContextPlugin_free_learn_GSHARE_COUNTER_0 + (1'b1 ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l123 = (((BranchContextPlugin_learn_BRANCH_FINAL_taken && BranchContextPlugin_free_learn_GSHARE_COUNTER_0[1]) && (! GSharePlugin_logic_onLearn_updated_0[1])) || (((! BranchContextPlugin_learn_BRANCH_FINAL_taken) && (! BranchContextPlugin_free_learn_GSHARE_COUNTER_0[1])) && GSharePlugin_logic_onLearn_updated_0[1]));
  assign GSharePlugin_logic_mem_write_valid = ((BranchContextPlugin_setup_learnValid && BranchContextPlugin_free_learn_Prediction_IS_BRANCH) && (! GSharePlugin_logic_onLearn_overflow));
  assign GSharePlugin_logic_mem_write_payload_address = GSharePlugin_logic_onLearn_hash;
  assign GSharePlugin_logic_mem_write_payload_data_0 = GSharePlugin_logic_onLearn_updated_0;
  assign DataCachePlugin_setup_writebackBusy = DataCachePlugin_logic_cache_io_writebackBusy;
  assign DataCachePlugin_setup_refillCompletions = DataCachePlugin_logic_cache_io_refillCompletions;
  assign DataCachePlugin_logic_load_hits = {Lsu2Plugin_setup_cacheLoad_cmd_valid,MmuPlugin_setup_cacheLoad_cmd_valid};
  assign DataCachePlugin_logic_load_hit = (|DataCachePlugin_logic_load_hits);
  assign _zz_DataCachePlugin_logic_load_hits_bools_0 = DataCachePlugin_logic_load_hits;
  assign DataCachePlugin_logic_load_hits_bools_0 = _zz_DataCachePlugin_logic_load_hits_bools_0[0];
  assign DataCachePlugin_logic_load_hits_bools_1 = _zz_DataCachePlugin_logic_load_hits_bools_0[1];
  always @(*) begin
    _zz_DataCachePlugin_logic_load_oh[0] = (DataCachePlugin_logic_load_hits_bools_0 && (! 1'b0));
    _zz_DataCachePlugin_logic_load_oh[1] = (DataCachePlugin_logic_load_hits_bools_1 && (! DataCachePlugin_logic_load_hits_bools_0));
  end

  assign DataCachePlugin_logic_load_oh = _zz_DataCachePlugin_logic_load_oh;
  assign _zz_DataCachePlugin_logic_load_ohHistory_0 = DataCachePlugin_logic_load_oh;
  assign DataCachePlugin_logic_load_ohHistory_0 = _zz_DataCachePlugin_logic_load_ohHistory_0;
  assign DataCachePlugin_logic_load_ohHistory_1 = _zz_DataCachePlugin_logic_load_ohHistory_1;
  assign DataCachePlugin_logic_load_ohHistory_2 = _zz_DataCachePlugin_logic_load_ohHistory_2;
  assign _zz_MmuPlugin_setup_cacheLoad_cmd_ready = DataCachePlugin_logic_load_oh[0];
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_virtual = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_virtual : Lsu2Plugin_setup_cacheLoad_cmd_payload_virtual);
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_size = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_size : Lsu2Plugin_setup_cacheLoad_cmd_payload_size);
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_redoOnDataHazard = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_redoOnDataHazard : Lsu2Plugin_setup_cacheLoad_cmd_payload_redoOnDataHazard);
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_unlocked = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_unlocked : Lsu2Plugin_setup_cacheLoad_cmd_payload_unlocked);
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_unique = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_unique : Lsu2Plugin_setup_cacheLoad_cmd_payload_unique);
  assign MmuPlugin_setup_cacheLoad_cmd_ready = _zz_MmuPlugin_setup_cacheLoad_cmd_ready;
  assign Lsu2Plugin_setup_cacheLoad_cmd_ready = DataCachePlugin_logic_load_oh[1];
  assign DataCachePlugin_logic_cache_io_load_cancels = (MmuPlugin_setup_cacheLoad_cancels | Lsu2Plugin_setup_cacheLoad_cancels);
  assign _zz_io_load_translated_physical = DataCachePlugin_logic_load_ohHistory_1[0];
  assign DataCachePlugin_logic_cache_io_load_translated_physical = (_zz_io_load_translated_physical ? MmuPlugin_setup_cacheLoad_translated_physical : Lsu2Plugin_setup_cacheLoad_translated_physical);
  assign DataCachePlugin_logic_cache_io_load_translated_abord = (_zz_io_load_translated_physical ? MmuPlugin_setup_cacheLoad_translated_abord : Lsu2Plugin_setup_cacheLoad_translated_abord);
  assign MmuPlugin_setup_cacheLoad_rsp_valid = (DataCachePlugin_logic_cache_io_load_rsp_valid && DataCachePlugin_logic_load_ohHistory_2[0]);
  assign MmuPlugin_setup_cacheLoad_rsp_payload_data = DataCachePlugin_logic_cache_io_load_rsp_payload_data;
  assign MmuPlugin_setup_cacheLoad_rsp_payload_fault = DataCachePlugin_logic_cache_io_load_rsp_payload_fault;
  assign MmuPlugin_setup_cacheLoad_rsp_payload_redo = DataCachePlugin_logic_cache_io_load_rsp_payload_redo;
  assign MmuPlugin_setup_cacheLoad_rsp_payload_refillSlot = DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlot;
  assign MmuPlugin_setup_cacheLoad_rsp_payload_refillSlotAny = DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlotAny;
  assign Lsu2Plugin_setup_cacheLoad_rsp_valid = (DataCachePlugin_logic_cache_io_load_rsp_valid && DataCachePlugin_logic_load_ohHistory_2[1]);
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_data = DataCachePlugin_logic_cache_io_load_rsp_payload_data;
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_fault = DataCachePlugin_logic_cache_io_load_rsp_payload_fault;
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_redo = DataCachePlugin_logic_cache_io_load_rsp_payload_redo;
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlot = DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlot;
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlotAny = DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlotAny;
  assign Lsu2Plugin_setup_cacheStore_cmd_ready = DataCachePlugin_logic_cache_io_store_cmd_ready;
  assign Lsu2Plugin_setup_cacheStore_rsp_valid = DataCachePlugin_logic_cache_io_store_rsp_valid;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_fault = DataCachePlugin_logic_cache_io_store_rsp_payload_fault;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_redo = DataCachePlugin_logic_cache_io_store_rsp_payload_redo;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlot = DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlot;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlotAny = DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlotAny;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_generationKo = DataCachePlugin_logic_cache_io_store_rsp_payload_generationKo;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_flush = DataCachePlugin_logic_cache_io_store_rsp_payload_flush;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_prefetch = DataCachePlugin_logic_cache_io_store_rsp_payload_prefetch;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_address = DataCachePlugin_logic_cache_io_store_rsp_payload_address;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_io = DataCachePlugin_logic_cache_io_store_rsp_payload_io;
  assign DataCachePlugin_mem_read_cmd_valid = DataCachePlugin_logic_cache_io_mem_read_cmd_valid;
  assign DataCachePlugin_mem_read_cmd_payload_id = DataCachePlugin_logic_cache_io_mem_read_cmd_payload_id;
  assign DataCachePlugin_mem_read_cmd_payload_address = DataCachePlugin_logic_cache_io_mem_read_cmd_payload_address;
  assign DataCachePlugin_mem_read_rsp_ready = DataCachePlugin_logic_cache_io_mem_read_rsp_ready;
  assign DataCachePlugin_mem_write_cmd_valid = DataCachePlugin_logic_cache_io_mem_write_cmd_valid;
  assign DataCachePlugin_mem_write_cmd_payload_last = DataCachePlugin_logic_cache_io_mem_write_cmd_payload_last;
  assign DataCachePlugin_mem_write_cmd_payload_fragment_address = DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_address;
  assign DataCachePlugin_mem_write_cmd_payload_fragment_data = DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_data;
  assign DataCachePlugin_mem_write_cmd_payload_fragment_id = DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_id;
  assign CommitPlugin_logic_ptr_commitRow = CommitPlugin_logic_ptr_commit;
  always @(*) begin
    CommitPlugin_logic_ptr_commitNext = CommitPlugin_logic_ptr_commit;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_logic_commit_lineCommited) begin
        CommitPlugin_logic_ptr_commitNext = (CommitPlugin_logic_ptr_commit + 5'h01);
      end
      if(CommitPlugin_logic_commit_rescheduleHit) begin
        CommitPlugin_logic_ptr_commitNext = CommitPlugin_logic_ptr_allocNext;
      end
    end
  end

  assign CommitPlugin_logic_ptr_full = ((CommitPlugin_logic_ptr_alloc ^ CommitPlugin_logic_ptr_free) == 5'h10);
  assign CommitPlugin_logic_ptr_canFree = (CommitPlugin_logic_ptr_free != CommitPlugin_logic_ptr_commit);
  assign CommitPlugin_setup_robLineMask_line = CommitPlugin_logic_ptr_commitNext[3:0];
  assign FrontendPlugin_allocated_ROB_ID = CommitPlugin_logic_ptr_alloc[3:0];
  assign FrontendPlugin_allocated_ROB_MSB_0 = CommitPlugin_logic_ptr_alloc[4];
  assign FrontendPlugin_allocated_haltRequest_CommitPlugin_l95 = CommitPlugin_logic_ptr_full;
  assign CommitPlugin_logic_ptr_allocNext = (CommitPlugin_logic_ptr_alloc + _zz_CommitPlugin_logic_ptr_allocNext);
  assign CommitPlugin_setup_isRobEmpty = CommitPlugin_logic_ptr_empty;
  assign CommitPlugin_logic_reschedule_commit_row = CommitPlugin_logic_reschedule_robId;
  assign CommitPlugin_logic_reschedule_commit_rowHit = (CommitPlugin_logic_reschedule_valid && (CommitPlugin_logic_reschedule_commit_row == _zz_CommitPlugin_logic_reschedule_commit_rowHit));
  assign CommitPlugin_logic_reschedule_age = (CommitPlugin_logic_reschedule_robId - _zz_CommitPlugin_logic_reschedule_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_0_age = (Lsu2Plugin_setup_sharedTrap_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_0_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_1_age = (Lsu2Plugin_setup_specialTrap_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_1_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_2_age = (EU0_BranchPlugin_setup_reschedule_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_2_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_3_age = (EnvCallPlugin_setup_reschedule_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_3_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_4_age = (EU0_CsrAccessPlugin_setup_trap_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_4_age);
  always @(*) begin
    CommitPlugin_logic_reschedule_portsLogic_hits[0] = (Lsu2Plugin_setup_sharedTrap_valid && (&{((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_4_age)),{((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_3_age)),{((! EU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_2_age)),{(_zz_CommitPlugin_logic_reschedule_portsLogic_hits || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_1),(_zz_CommitPlugin_logic_reschedule_portsLogic_hits_2 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_3)}}}}));
    CommitPlugin_logic_reschedule_portsLogic_hits[1] = (Lsu2Plugin_setup_specialTrap_valid && (&{((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_4_age)),{((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_3_age)),{((! EU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_2_age)),{(_zz_CommitPlugin_logic_reschedule_portsLogic_hits_4 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_5),(_zz_CommitPlugin_logic_reschedule_portsLogic_hits_6 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_7)}}}}));
    CommitPlugin_logic_reschedule_portsLogic_hits[2] = (EU0_BranchPlugin_setup_reschedule_valid && (&{((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_4_age)),{((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_3_age)),{((! Lsu2Plugin_setup_specialTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age < CommitPlugin_logic_reschedule_portsLogic_perPort_1_age)),{((! Lsu2Plugin_setup_sharedTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age)),((! CommitPlugin_logic_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age < CommitPlugin_logic_reschedule_age))}}}}));
    CommitPlugin_logic_reschedule_portsLogic_hits[3] = (EnvCallPlugin_setup_reschedule_valid && (&{((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_4_age)),{((! EU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age < CommitPlugin_logic_reschedule_portsLogic_perPort_2_age)),{((! Lsu2Plugin_setup_specialTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age < CommitPlugin_logic_reschedule_portsLogic_perPort_1_age)),{(_zz_CommitPlugin_logic_reschedule_portsLogic_hits_8 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_9),(_zz_CommitPlugin_logic_reschedule_portsLogic_hits_10 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_11)}}}}));
    CommitPlugin_logic_reschedule_portsLogic_hits[4] = (EU0_CsrAccessPlugin_setup_trap_valid && (&{((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_portsLogic_perPort_3_age)),{((! EU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_portsLogic_perPort_2_age)),{((! Lsu2Plugin_setup_specialTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_portsLogic_perPort_1_age)),{((! Lsu2Plugin_setup_sharedTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age)),((! CommitPlugin_logic_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_age))}}}}));
  end

  assign when_CommitPlugin_l131 = (|CommitPlugin_logic_reschedule_portsLogic_hits);
  assign _zz_CommitPlugin_logic_reschedule_trap = CommitPlugin_logic_reschedule_portsLogic_hits[0];
  assign _zz_CommitPlugin_logic_reschedule_trap_1 = CommitPlugin_logic_reschedule_portsLogic_hits[1];
  assign _zz_CommitPlugin_logic_reschedule_trap_2 = CommitPlugin_logic_reschedule_portsLogic_hits[2];
  assign _zz_CommitPlugin_logic_reschedule_trap_3 = CommitPlugin_logic_reschedule_portsLogic_hits[3];
  assign _zz_CommitPlugin_logic_reschedule_trap_4 = CommitPlugin_logic_reschedule_portsLogic_hits[4];
  assign CommitPlugin_setup_jump_valid = (CommitPlugin_logic_reschedule_fresh && (! CommitPlugin_logic_reschedule_trap));
  assign CommitPlugin_setup_jump_payload_pc = CommitPlugin_logic_reschedule_pcTarget;
  assign CommitPlugin_logic_reschedule_reschedulePort_valid = CommitPlugin_logic_reschedule_fresh;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_robId = CommitPlugin_logic_reschedule_robId;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_trap = CommitPlugin_logic_reschedule_trap;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_cause = CommitPlugin_logic_reschedule_cause;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_tval = CommitPlugin_logic_reschedule_tval;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_reason = CommitPlugin_logic_reschedule_reason;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_skipCommit = CommitPlugin_logic_reschedule_skipCommit;
  always @(*) begin
    CommitPlugin_logic_commit_rescheduleHit = 1'b0;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_0_enable) begin
        if(CommitPlugin_logic_commit_continue) begin
          if(when_CommitPlugin_l207) begin
            CommitPlugin_logic_commit_rescheduleHit = 1'b1;
          end
        end
      end
    end
  end

  assign CommitPlugin_logic_commit_active = _zz_CommitPlugin_logic_commit_active_1[0];
  always @(*) begin
    CommitPlugin_logic_commit_maskComb = CommitPlugin_logic_commit_mask;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_0_enable) begin
        if(CommitPlugin_logic_commit_continue) begin
          if(when_CommitPlugin_l203) begin
            CommitPlugin_logic_commit_maskComb[0] = 1'b0;
          end
        end
      end
    end
  end

  assign CommitPlugin_logic_commit_lineCommited = ((CommitPlugin_logic_commit_maskComb & CommitPlugin_logic_commit_active) == 1'b0);
  always @(*) begin
    CommitPlugin_logic_commit_event_mask = 1'b0;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_0_enable) begin
        if(CommitPlugin_logic_commit_continue) begin
          if(when_CommitPlugin_l203) begin
            CommitPlugin_logic_commit_event_mask[0] = 1'b1;
          end
        end
      end
    end
  end

  assign CommitPlugin_logic_commit_event_robId = CommitPlugin_logic_ptr_commit[3:0];
  always @(*) begin
    CommitPlugin_logic_commit_lineEvent_valid = 1'b0;
    if(when_CommitPlugin_l194) begin
      if(when_CommitPlugin_l217) begin
        CommitPlugin_logic_commit_lineEvent_valid = 1'b1;
      end
    end
  end

  assign CommitPlugin_logic_commit_lineEvent_payload_mask = (CommitPlugin_logic_commit_active ^ CommitPlugin_logic_commit_maskComb);
  assign CommitPlugin_logic_commit_lineEvent_payload_robId = CommitPlugin_logic_ptr_commit[3:0];
  assign CommitPlugin_logic_commit_reschedulePort_valid = CommitPlugin_logic_commit_rescheduleHit;
  assign CommitPlugin_logic_commit_reschedulePort_payload_robId = CommitPlugin_logic_reschedule_robId;
  assign CommitPlugin_logic_commit_reschedulePort_payload_robIdNext = CommitPlugin_logic_ptr_allocNext[3:0];
  assign CommitPlugin_logic_commit_reschedulePort_payload_trap = CommitPlugin_logic_reschedule_trap;
  assign CommitPlugin_logic_commit_reschedulePort_payload_cause = CommitPlugin_logic_reschedule_cause;
  assign CommitPlugin_logic_commit_reschedulePort_payload_tval = CommitPlugin_logic_reschedule_tval;
  assign CommitPlugin_logic_commit_reschedulePort_payload_reason = CommitPlugin_logic_reschedule_reason;
  assign CommitPlugin_logic_commit_reschedulePort_payload_skipCommit = CommitPlugin_logic_reschedule_skipCommit;
  always @(*) begin
    CommitPlugin_logic_commit_headNext = CommitPlugin_logic_commit_head;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_logic_commit_rescheduleHit) begin
        CommitPlugin_logic_commit_headNext = CommitPlugin_logic_ptr_allocNext[3:0];
      end
    end
  end

  assign CommitPlugin_logic_commit_head = _zz_CommitPlugin_logic_commit_head[3:0];
  assign CommitPlugin_logic_commit_continue = 1'b1;
  assign when_CommitPlugin_l194 = (! CommitPlugin_logic_ptr_empty);
  assign CommitPlugin_commit_slot_0_enable = (CommitPlugin_logic_commit_mask[0] && CommitPlugin_logic_commit_active[0]);
  assign CommitPlugin_commit_slot_0_readyForCommit = CommitPlugin_logic_ptr_robLineMaskRsp[0];
  assign CommitPlugin_commit_slot_0_rescheduleHitSlot = (CommitPlugin_logic_reschedule_commit_rowHit && 1'b1);
  assign when_CommitPlugin_l203 = (CommitPlugin_commit_slot_0_readyForCommit && (! (CommitPlugin_commit_slot_0_rescheduleHitSlot && CommitPlugin_logic_reschedule_skipCommit)));
  assign when_CommitPlugin_l207 = (CommitPlugin_commit_slot_0_rescheduleHitSlot && (CommitPlugin_logic_reschedule_skipCommit || CommitPlugin_commit_slot_0_readyForCommit));
  assign when_CommitPlugin_l211 = ((! CommitPlugin_commit_slot_0_readyForCommit) || CommitPlugin_commit_slot_0_rescheduleHitSlot);
  assign when_CommitPlugin_l217 = (CommitPlugin_logic_commit_lineCommited || CommitPlugin_logic_commit_rescheduleHit);
  assign CommitPlugin_logic_free_lineEventStream_valid = CommitPlugin_logic_commit_lineEvent_valid;
  assign CommitPlugin_logic_free_lineEventStream_payload_robId = CommitPlugin_logic_commit_lineEvent_payload_robId;
  assign CommitPlugin_logic_free_lineEventStream_payload_mask = CommitPlugin_logic_commit_lineEvent_payload_mask;
  assign CommitPlugin_logic_free_lineEventStream_ready = CommitPlugin_logic_free_lineEventStream_fifo_io_push_ready;
  assign CommitPlugin_logic_free_robHit = (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_robId == _zz_CommitPlugin_logic_free_robHit);
  assign CommitPlugin_logic_free_hit = (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_valid && CommitPlugin_logic_free_robHit);
  assign CommitPlugin_logic_free_lineEventStream_fifo_io_pop_ready = (CommitPlugin_logic_free_robHit && CommitPlugin_logic_ptr_canFree);
  assign CommitPlugin_logic_free_port_valid = CommitPlugin_logic_ptr_canFree;
  assign CommitPlugin_logic_free_port_payload_robId = CommitPlugin_logic_ptr_free[3:0];
  assign CommitPlugin_logic_free_port_payload_commited = (CommitPlugin_logic_free_hit ? CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_mask : 1'b0);
  assign robToPc_valid = FrontendPlugin_allocated_isFireing;
  assign robToPc_robId = FrontendPlugin_allocated_ROB_ID;
  assign robToPc_pc_0 = FrontendPlugin_allocated_PC_0;
  assign commit_robId = CommitPlugin_logic_commit_event_robId;
  assign commit_mask = CommitPlugin_logic_commit_event_mask;
  assign reschedule_valid = CommitPlugin_logic_commit_reschedulePort_valid;
  assign reschedule_payload_robId = CommitPlugin_logic_commit_reschedulePort_payload_robId;
  assign reschedule_payload_robIdNext = CommitPlugin_logic_commit_reschedulePort_payload_robIdNext;
  assign reschedule_payload_trap = CommitPlugin_logic_commit_reschedulePort_payload_trap;
  assign reschedule_payload_cause = CommitPlugin_logic_commit_reschedulePort_payload_cause;
  assign reschedule_payload_tval = CommitPlugin_logic_commit_reschedulePort_payload_tval;
  assign reschedule_payload_reason = CommitPlugin_logic_commit_reschedulePort_payload_reason;
  assign reschedule_payload_skipCommit = CommitPlugin_logic_commit_reschedulePort_payload_skipCommit;
  assign rescheduleReason = CommitPlugin_logic_reschedule_reason;
  assign commit_pc_0 = _zz_commit_pc_0_1[31 : 0];
  assign CommitDebugFilterPlugin_logic_commits = ({16'd0,_zz_CommitDebugFilterPlugin_logic_commits} <<< 5'd16);
  assign PrivilegedPlugin_logic_defaultTrap_csrPrivilege = EU0_CsrAccessPlugin_setup_onDecodeAddress[9 : 8];
  assign PrivilegedPlugin_logic_defaultTrap_csrReadOnly = (&EU0_CsrAccessPlugin_setup_onDecodeAddress[11 : 10]);
  assign when_PrivilegedPlugin_l165 = ((PrivilegedPlugin_logic_defaultTrap_csrReadOnly && EU0_CsrAccessPlugin_setup_onDecodeWrite) || (PrivilegedPlugin_setup_privilege < PrivilegedPlugin_logic_defaultTrap_csrPrivilege));
  always @(*) begin
    PrivilegedPlugin_logic_machine_mstatus_sd = 1'b0;
    if(when_PrivilegedPlugin_l393) begin
      PrivilegedPlugin_logic_machine_mstatus_sd = 1'b1;
    end
  end

  assign when_PrivilegedPlugin_l393 = (PrivilegedPlugin_logic_machine_mstatus_fs == 2'b11);
  assign PrivilegedPlugin_logic_supervisor_sip_seipOr = (PrivilegedPlugin_logic_supervisor_sip_seipSoft || PrivilegedPlugin_logic_supervisor_sip_seipInput);
  assign PrivilegedPlugin_logic_supervisor_sip_seipMasked = (PrivilegedPlugin_logic_supervisor_sip_seipOr && PrivilegedPlugin_logic_machine_mideleg_se);
  assign PrivilegedPlugin_logic_supervisor_sip_stipMasked = (PrivilegedPlugin_logic_supervisor_sip_stip && PrivilegedPlugin_logic_machine_mideleg_st);
  assign PrivilegedPlugin_logic_supervisor_sip_ssipMasked = (PrivilegedPlugin_logic_supervisor_sip_ssip && PrivilegedPlugin_logic_machine_mideleg_ss);
  assign _zz_when_PrivilegedPlugin_l644 = (PrivilegedPlugin_logic_supervisor_sip_ssip && PrivilegedPlugin_logic_supervisor_sie_ssie);
  assign _zz_when_PrivilegedPlugin_l644_1 = (PrivilegedPlugin_logic_supervisor_sip_stip && PrivilegedPlugin_logic_supervisor_sie_stie);
  assign _zz_when_PrivilegedPlugin_l644_2 = (PrivilegedPlugin_logic_supervisor_sip_seipOr && PrivilegedPlugin_logic_supervisor_sie_seie);
  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_ready = PrivilegedPlugin_logic_reschedule_ready;
    if(when_Stream_l369) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_ready = 1'b1;
    end
  end

  assign when_Stream_l369 = (! PrivilegedPlugin_logic_reschedule_valid);
  assign PrivilegedPlugin_logic_reschedule_valid = PrivilegedPlugin_logic_rescheduleUnbuffered_rValid;
  assign PrivilegedPlugin_logic_reschedule_payload_cause = PrivilegedPlugin_logic_rescheduleUnbuffered_rData_cause;
  assign PrivilegedPlugin_logic_reschedule_payload_epc = PrivilegedPlugin_logic_rescheduleUnbuffered_rData_epc;
  assign PrivilegedPlugin_logic_reschedule_payload_tval = PrivilegedPlugin_logic_rescheduleUnbuffered_rData_tval;
  assign PrivilegedPlugin_logic_reschedule_payload_fromCommit = PrivilegedPlugin_logic_rescheduleUnbuffered_rData_fromCommit;
  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_valid = (CommitPlugin_logic_commit_reschedulePort_valid && CommitPlugin_logic_commit_reschedulePort_payload_trap);
    if(when_PrivilegedPlugin_l592) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_valid = 1'b1;
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_payload_cause = CommitPlugin_logic_commit_reschedulePort_payload_cause;
    if(when_PrivilegedPlugin_l592) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_payload_cause = DecoderPlugin_setup_exceptionPort_payload_cause;
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc = _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_1[31 : 0];
    if(when_PrivilegedPlugin_l592) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc = DecoderPlugin_setup_exceptionPort_payload_epc;
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_payload_tval = CommitPlugin_logic_commit_reschedulePort_payload_tval;
    if(when_PrivilegedPlugin_l592) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_payload_tval = DecoderPlugin_setup_exceptionPort_payload_tval;
    end
  end

  assign PrivilegedPlugin_logic_rescheduleUnbuffered_payload_fromCommit = (CommitPlugin_logic_commit_reschedulePort_valid && CommitPlugin_logic_commit_reschedulePort_payload_trap);
  assign when_PrivilegedPlugin_l592 = (DecoderPlugin_setup_exceptionPort_valid && (! PrivilegedPlugin_logic_rescheduleUnbuffered_payload_fromCommit));
  assign PrivilegedPlugin_logic_targetMachine = 1'b1;
  always @(*) begin
    PrivilegedPlugin_logic_reschedule_ready = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
        PrivilegedPlugin_logic_reschedule_ready = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  assign ALU0_IntFormatPlugin_logic_stages_0_hits = {ALU0_ShiftPlugin_setup_intFormatPort_valid,ALU0_IntAluPlugin_setup_intFormatPort_valid};
  assign ALU0_IntFormatPlugin_logic_stages_0_wb_valid = (ALU0_ExecutionUnitBase_pipeline_execute_0_valid && (|ALU0_IntFormatPlugin_logic_stages_0_hits));
  assign ALU0_IntFormatPlugin_logic_stages_0_raw = ((ALU0_IntFormatPlugin_logic_stages_0_hits[0] ? ALU0_IntAluPlugin_setup_intFormatPort_payload : 32'h00000000) | (ALU0_IntFormatPlugin_logic_stages_0_hits[1] ? ALU0_ShiftPlugin_setup_intFormatPort_payload : 32'h00000000));
  assign ALU0_IntFormatPlugin_logic_stages_0_wb_payload = ALU0_IntFormatPlugin_logic_stages_0_raw;
  always @(*) begin
    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL)
      1'b0 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
      end
      default : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = {ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 12],12'h000};
      end
    endcase
  end

  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  always @(*) begin
    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL)
      2'b00 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
      end
      2'b01 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {{20{_zz__zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2[11]}}, _zz__zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2};
      end
      2'b10 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU0_ExecutionUnitBase_pipeline_fetch_0_PC;
      end
      default : begin
      end
    endcase
  end

  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  always @(*) begin
    ALU0_SrcPlugin_logic_addsub_rs2Patched = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
    if(ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT) begin
      ALU0_SrcPlugin_logic_addsub_rs2Patched = (~ ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
    end
    if(ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO) begin
      ALU0_SrcPlugin_logic_addsub_rs2Patched = 32'h00000000;
    end
  end

  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(_zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB) + $signed(_zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1));
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS = ((ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31] == ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31]) ? ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB[31] : (ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED ? ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31] : ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]));
  assign ALU0_IntAluPlugin_setup_intFormatPort_valid = ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL;
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        ALU0_IntAluPlugin_logic_process_bitwise = (ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 & ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        ALU0_IntAluPlugin_logic_process_bitwise = (ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 | ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
      default : begin
        ALU0_IntAluPlugin_logic_process_bitwise = (ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 ^ ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
    endcase
  end

  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_BITWISE : begin
        ALU0_IntAluPlugin_logic_process_result = ALU0_IntAluPlugin_logic_process_bitwise;
      end
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : begin
        ALU0_IntAluPlugin_logic_process_result = _zz_ALU0_IntAluPlugin_logic_process_result;
      end
      default : begin
        ALU0_IntAluPlugin_logic_process_result = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
      end
    endcase
  end

  assign ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT = ALU0_IntAluPlugin_logic_process_result;
  assign ALU0_IntAluPlugin_setup_intFormatPort_payload = ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT;
  assign ALU0_ShiftPlugin_setup_intFormatPort_valid = ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL;
  assign ALU0_ShiftPlugin_logic_process_amplitude = _zz_ALU0_ShiftPlugin_logic_process_amplitude;
  assign ALU0_ShiftPlugin_logic_process_reversed = (ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT ? _zz_ALU0_ShiftPlugin_logic_process_reversed : ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1);
  assign ALU0_ShiftPlugin_logic_process_shifted = _zz_ALU0_ShiftPlugin_logic_process_shifted[31:0];
  assign ALU0_ShiftPlugin_logic_process_patched = (ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT ? _zz_ALU0_ShiftPlugin_logic_process_patched : ALU0_ShiftPlugin_logic_process_shifted);
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT = ALU0_ShiftPlugin_logic_process_patched;
  assign ALU0_ShiftPlugin_setup_intFormatPort_payload = ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT;
  assign EU0_IntFormatPlugin_logic_stages_0_hits = {EU0_CsrAccessPlugin_setup_intFormatPort_valid,{EU0_BranchPlugin_setup_intFormatPort_valid,{EU0_DivPlugin_setup_intFormatPort_valid,EU0_MulPlugin_setup_intFormatPort_valid}}};
  assign EU0_IntFormatPlugin_logic_stages_0_wb_valid = (EU0_ExecutionUnitBase_pipeline_execute_2_valid && (|EU0_IntFormatPlugin_logic_stages_0_hits));
  assign EU0_IntFormatPlugin_logic_stages_0_raw = (((EU0_IntFormatPlugin_logic_stages_0_hits[0] ? EU0_MulPlugin_setup_intFormatPort_payload : 32'h00000000) | (EU0_IntFormatPlugin_logic_stages_0_hits[1] ? EU0_DivPlugin_setup_intFormatPort_payload : 32'h00000000)) | ((EU0_IntFormatPlugin_logic_stages_0_hits[2] ? EU0_BranchPlugin_setup_intFormatPort_payload : 32'h00000000) | (EU0_IntFormatPlugin_logic_stages_0_hits[3] ? EU0_CsrAccessPlugin_setup_intFormatPort_payload : 32'h00000000)));
  assign EU0_IntFormatPlugin_logic_stages_0_wb_payload = EU0_IntFormatPlugin_logic_stages_0_raw;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
  end

  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(EU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL)
      2'b00 : begin
        _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
      end
      2'b01 : begin
        _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {{20{_zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2[11]}}, _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2};
      end
      2'b10 : begin
        _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {{20{_zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2_1[11]}}, _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2_1};
      end
      default : begin
      end
    endcase
  end

  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  always @(*) begin
    EU0_SrcPlugin_logic_addsub_rs2Patched = EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
    if(EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT) begin
      EU0_SrcPlugin_logic_addsub_rs2Patched = (~ EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO) begin
      EU0_SrcPlugin_logic_addsub_rs2Patched = 32'h00000000;
    end
  end

  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB) + $signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1));
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS = ((EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31] == EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31]) ? EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB[31] : (EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED ? EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31] : EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]));
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED = EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED = EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT = (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_SIGNED && EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED[31]);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT = (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED && EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED[31]);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED = ((EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT ? (~ EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED) : EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED) + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED = ((EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT ? (~ EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED) : EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED) + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED);
  assign EU0_MulPlugin_setup_intFormatPort_valid = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL;
  assign EU0_MulPlugin_logic_wake_wakeRobsSel = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL;
  assign EU0_MulPlugin_logic_wake_wakeRegFileSel = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1 = {(EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_SIGNED && EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1[31]),EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1};
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2 = {(EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED && EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2[31]),EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2};
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_0 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[0] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[1] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[2] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_5 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[3] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_7 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[4] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_9 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[5] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_11 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[6] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_13 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[7] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_15 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[8] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_17 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[9] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_19 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[10] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_21 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[11] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_23 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[12] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_25 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[13] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_27 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[14] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_29 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[15] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_31 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[16] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_33 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[17] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_35 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[18] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_37 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[19] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_39 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[20] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_41 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[21] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_43 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[22] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_45 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[23] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_47 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[24] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_49 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[25] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_51 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[26] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_53 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[27] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_55 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[28] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_57 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[29] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_59 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[30] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_61 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[31] ? EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[31 : 0] : 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_63 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_63;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0[20 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_0[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_1 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_1[20 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_2 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_2[20 : 2] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_3 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_3[20 : 3] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_5[17 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1[20 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_7[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_1 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_1[20 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_9[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_2 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_2[20 : 2] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_11[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_3 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_3[20 : 3] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_13[17 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2[20 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_15[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_1 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_1[20 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_17[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_2 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_2[20 : 2] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_19[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_3 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_3[20 : 3] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_21[17 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3[20 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_23[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_1 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_1[20 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_25[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_2 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_2[20 : 2] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_27[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_3 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_3[20 : 3] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_29[17 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4[20 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_31[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_1 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_1[20 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_33[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_2 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_2[20 : 2] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_35[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_3 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_3[20 : 3] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_37[17 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5[20 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_39[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_1 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_1[20 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_41[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_2 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_2[11 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_0[31 : 21];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_2[20 : 12] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2[8 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_3 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_3[12 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1[31 : 20];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_3[20 : 13] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4[7 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3[31 : 19];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6[19 : 13] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6[6 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_1 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_1[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_5[31 : 18];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_1[19 : 14] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8[5 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_2 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_2[19 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_43[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_3 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_3[19 : 2] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_45[17 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7[20 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_47[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_1 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_1[20 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_49[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_2 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_2[11 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_7[31 : 21];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_2[20 : 12] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10[8 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_3 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_3[12 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_9[31 : 20];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_3[20 : 13] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12[7 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_11[31 : 19];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8[19 : 13] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14[6 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_1 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_1[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_13[31 : 18];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_1[19 : 14] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16[5 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_2 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_2[19 : 1] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_51[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_3 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_3[19 : 2] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_53[17 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_9 = 32'h00000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_9[31 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_55[31 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_10 = 32'h00000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_10[31 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_57[31 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_11 = 11'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_11[10 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_15[31 : 21];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_12 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_12[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_17[31 : 20];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_13 = 13'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_13[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_19[31 : 19];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_14 = 14'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_14[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_21[31 : 18];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_15 = 32'h00000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_15[31 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_59[31 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_16 = 32'h00000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_16[31 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_61[31 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_17 = 32'h00000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_17[31 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_64[31 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_18 = 11'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_18[10 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_23[31 : 21];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_19 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_19[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_25[31 : 20];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_20 = 13'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_20[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_27[31 : 19];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_21 = 14'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_21[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_29[31 : 18];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_22 = 11'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_22[10 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_31[31 : 21];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_23 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_23[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_33[31 : 20];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_24 = 13'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_24[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_35[31 : 19];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_25 = 14'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_25[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_37[31 : 18];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_26 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_26[23 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_18[23 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_27 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_27[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_20[22 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_28 = 11'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_28[10 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_39[31 : 21];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_29 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_29[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_41[31 : 20];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_30 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_30[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2[31 : 9];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_31 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_31[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_4[30 : 8];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_32 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_32[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_6[29 : 7];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_33 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_33[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_8[28 : 6];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_34 = 13'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_34[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_43[31 : 19];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_35 = 14'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_35[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_45[31 : 18];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_36 = 22'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_36[21 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_22[21 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_37 = 21'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_37[20 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_24[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_38 = 20'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_38[19 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_26[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_39 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_39[18 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_28[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_40 = 11'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_40[10 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_47[31 : 21];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_41 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_41[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_49[31 : 20];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_42 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_42[18 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_10[27 : 9];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_43 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_43[18 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_12[26 : 8];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_44 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_44[18 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_14[25 : 7];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_45 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_45[18 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_16[24 : 6];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_46 = 13'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_46[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_51[31 : 19];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_47 = 14'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_47[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_53[31 : 18];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_48 = 18'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_48[17 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_30[17 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_49 = 17'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_49[16 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_32[16 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_50 = 16'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_50[15 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_34[15 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_51 = 15'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_51[14 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_36[14 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_52 = 14'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_52[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_38[13 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_53 = 13'h0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_53[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_40[12 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_54 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_54[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_42[11 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_55 = 11'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_55[10 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_44[10 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_56 = 10'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_56[9 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_46[9 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_57 = 9'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_57[8 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_48[8 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_58 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_58[7 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_50[7 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_59 = 7'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_59[6 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_52[6 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_60 = 6'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_60[5 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_54[5 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_61 = 5'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_61[4 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_56[4 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_62 = 4'b0000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_62[3 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_58[3 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_63 = 3'b000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_63[2 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_60[2 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_64 = 2'b00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_64[1 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_62[1 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_65 = 1'b0;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_65[0 : 0] = EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_63[0 : 0];
  end

  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8_7);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_9 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_9;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_10 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_10;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_11 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_11;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_12 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_12;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_13 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_13;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_14 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_14;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_15 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_15;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_16 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_16;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_17 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_17;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_18 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_18;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_19 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_19;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_20 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_20;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_21 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_21;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_22 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_22;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_23 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_23;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_24 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_24;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_25 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_25;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_26 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_26;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_27 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_27;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_28 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_28;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_29 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_29;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_30 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_30;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_31 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_31;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_32 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_32;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_33 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_33;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_34 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_34;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_35 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_35;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_36 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_36;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_37 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_37;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_38 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_38;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_39 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_39;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_40 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_40;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_41 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_41;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_42 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_42;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_43 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_43;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_44 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_44;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_45 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_45;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_46 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_46;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_47 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_47;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_48 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_48;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_49 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_49;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_50 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_50;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_51 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_51;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_52 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_52;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_53 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_53;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_54 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_54;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_55 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_55;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_56 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_56;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_57 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_57;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_58 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_58;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_59 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_59;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_60 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_60;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_61 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_61;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_62 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_62;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_63 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_63;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_64 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_64;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_65 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_65;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0 = 28'h0000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0[22 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0[27 : 24] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_7[3 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_1 = 28'h0000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_1[26 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1[22 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_2 = 28'h0000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_2[27 : 8] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_2[19 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_3 = 28'h0000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_3[27 : 12] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_3[15 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_4 = 28'h0000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_4[27 : 16] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_4[11 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_5 = 28'h0000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_5[27 : 20] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_5[7 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_6 = 28'h0000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_6[27 : 21] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_6[6 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_7 = 28'h0000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_7[27 : 25] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_8[2 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1[23 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_9[23 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_1 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_1[18 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_7[22 : 4];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_1[23 : 19] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_49[4 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_2 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_2[2 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_2[22 : 20];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_2[23 : 3] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_16[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_3 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_3[6 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_3[22 : 16];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_3[19 : 9] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_22[10 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_3[23 : 20] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_50[3 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_4 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_4[10 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_4[22 : 12];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_4[23 : 12] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_26[11 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_5 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_5[14 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_5[22 : 8];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_5[23 : 15] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_37[8 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_6 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_6[14 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_6[21 : 7];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_6[23 : 16] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_38[7 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_7 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_7[18 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_8[21 : 3];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_7[23 : 21] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_51[2 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2[23 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_10[23 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_1 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_1[10 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_11[10 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_1[23 : 12] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_27[11 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_2 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_2[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_12[11 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_2[22 : 12] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_28[10 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_2[23 : 23] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_54[0 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_3 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_3[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_13[12 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_3[23 : 13] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_36[10 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_4 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_4[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_14[13 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_4[23 : 16] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_39[7 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_5 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_5[23 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_15[22 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_6 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_6[23 : 3] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_17[20 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_7 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_7[14 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_18[10 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_7[23 : 16] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_40[7 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_19[11 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3[23 : 12] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_41[11 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_1 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_1[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_20[12 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_1[23 : 13] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_48[10 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_2 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_2[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_21[13 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_2[23 : 17] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_52[6 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_3 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_3[15 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_23[11 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_3[23 : 18] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_53[5 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_4 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_4[16 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_24[12 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_4[23 : 19] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_9[28 : 24];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_5 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_5[17 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_25[13 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_5[23 : 19] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_49[9 : 5];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_6 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_6[19 : 8] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_29[11 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_6[23 : 20] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_55[3 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_7 = 24'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_7[23 : 8] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_30[15 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_31[22 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_1 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_1[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_32[22 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_2 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_2[22 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_33[22 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_3 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_3[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_34[12 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_3[22 : 13] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_56[9 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_4 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_4[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_35[13 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_4[22 : 14] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_57[8 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_5 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_5[22 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_42[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_6 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_6[22 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_43[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_7 = 23'h000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_7[22 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_44[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5[18 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_45[18 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_1 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_1[12 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_46[12 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_1[18 : 13] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_60[5 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_2 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_2[13 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_47[13 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_2[18 : 14] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_61[4 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_3 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_3[17 : 7] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_16[31 : 21];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_3[18 : 18] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_65[0 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_4 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_4[18 : 7] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_50[15 : 4];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_5 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_5[18 : 7] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_26[23 : 12];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_6 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_6[18 : 7] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_37[20 : 9];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_7 = 19'h00000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_7[18 : 7] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_38[19 : 8];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6[11 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_51[14 : 3];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_1 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_1[8 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_10[31 : 24];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_1[11 : 9] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_63[2 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_2 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_2[11 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_27[22 : 12];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_3 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_3[11 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_54[11 : 1];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_4 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_4[11 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_36[21 : 11];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_5 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_5[11 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_39[18 : 8];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_6 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_6[9 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_15[31 : 23];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_6[11 : 10] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_64[1 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_7 = 12'h000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_7[11 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_17[31 : 21];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_7 = 3'b000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_7[2 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_40[10 : 8];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8[7 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_58[7 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_1 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_1[7 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_59[6 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_2 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_2[7 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_48[17 : 11];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_3 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_3[7 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_52[13 : 7];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_4 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_4[7 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_53[12 : 6];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_5 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_5[3 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_9[31 : 29];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_5[7 : 4] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_62[3 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_6 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_6[7 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_49[16 : 10];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_7 = 8'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_7[7 : 1] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_55[10 : 4];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_9 = 7'h00;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_9[6 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_30[22 : 16];
  end

  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0_15);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1_15);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2_15);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3_15);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4_15);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5_15);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6_15);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_7 = _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_7;
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_8 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8_15);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_9 = _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_9;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0 = 67'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0[30 : 0] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0[30 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0[59 : 33] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_3[26 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_1 = 67'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_1[54 : 28] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_1[26 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_1[66 : 56] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_8[10 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_2 = 67'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_2[55 : 29] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_2[26 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_2[63 : 57] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_9[6 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_3 = 67'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_3[66 : 41] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_4[25 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_4 = 67'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_4[66 : 45] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_5[21 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_5 = 67'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_5[66 : 52] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_6[14 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_6 = 67'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_6[55 : 53] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_7[2 : 0];
  end

  assign EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_7 + _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0_14);
  assign EU0_MulPlugin_setup_intFormatPort_payload = (EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_HIGH ? EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0[63 : 32] : EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_2_adders_0[31 : 0]);
  assign EU0_DivPlugin_setup_intFormatPort_valid = EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL;
  assign EU0_DivPlugin_logic_wake_wakeRobsSel = EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL;
  assign EU0_DivPlugin_logic_wake_wakeRegFileSel = EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_DIV_REVERT_RESULT = ((EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT ^ (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT && (! EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM))) && (! (((EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED == 32'h00000000) && EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED) && (! EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM))));
  assign toplevel_EU0_DivPlugin_logic_div_io_cmd_fire = (EU0_DivPlugin_logic_div_io_cmd_valid && EU0_DivPlugin_logic_div_io_cmd_ready);
  assign when_DivPlugin_l76 = (EU0_ExecutionUnitBase_pipeline_execute_0_ready || EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed);
  assign EU0_DivPlugin_logic_div_io_cmd_valid = ((EU0_ExecutionUnitBase_pipeline_execute_0_valid && EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL) && (! EU0_DivPlugin_logic_feed_cmdSent));
  assign EU0_ExecutionUnitBase_pipeline_execute_0_haltRequest_DivPlugin_l83 = ((EU0_ExecutionUnitBase_pipeline_execute_0_valid && EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL) && (! EU0_DivPlugin_logic_feed_cmdSent));
  assign EU0_ExecutionUnitBase_pipeline_execute_1_haltRequest_DivPlugin_l91 = ((EU0_ExecutionUnitBase_pipeline_execute_1_valid && EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_SEL) && (! EU0_DivPlugin_logic_div_io_rsp_valid));
  assign EU0_DivPlugin_logic_rsp_selected = (EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_REM ? _zz_EU0_DivPlugin_logic_rsp_selected : EU0_DivPlugin_logic_div_io_rsp_payload_result);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT = EU0_DivPlugin_logic_rsp_selected;
  assign EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT = _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_1[31:0];
  assign EU0_DivPlugin_setup_intFormatPort_payload = EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_DIV_RESULT;
  assign EU0_BranchPlugin_setup_intFormatPort_valid = EU0_ExecutionUnitBase_pipeline_execute_2_BranchPlugin_SEL;
  assign EU0_BranchPlugin_logic_wake_wakeRobsSel = EU0_ExecutionUnitBase_pipeline_execute_2_BranchPlugin_SEL;
  assign EU0_BranchPlugin_logic_wake_wakeRegFileSel = EU0_ExecutionUnitBase_pipeline_execute_2_BranchPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ = ($signed(EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1) == $signed(EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2));
  assign switch_Misc_l241 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[14 : 12];
  always @(*) begin
    casez(switch_Misc_l241)
      3'b000 : begin
        _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ;
      end
      3'b001 : begin
        _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = (! EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ);
      end
      3'b1?1 : begin
        _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = (! EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS);
      end
      default : begin
        _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
      end
    endcase
  end

  always @(*) begin
    case(EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = 1'b1;
      end
      default : begin
        _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
      end
    endcase
  end

  assign EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1;
  always @(*) begin
    case(EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        EU0_BranchPlugin_logic_process_target_a = EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1;
      end
      default : begin
        EU0_BranchPlugin_logic_process_target_a = EU0_ExecutionUnitBase_pipeline_execute_0_PC;
      end
    endcase
  end

  always @(*) begin
    case(EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        EU0_BranchPlugin_logic_process_target_b = {{11{_zz_EU0_BranchPlugin_logic_process_target_b[20]}}, _zz_EU0_BranchPlugin_logic_process_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        EU0_BranchPlugin_logic_process_target_b = {{20{_zz_EU0_BranchPlugin_logic_process_target_b_1[11]}}, _zz_EU0_BranchPlugin_logic_process_target_b_1};
      end
      default : begin
        EU0_BranchPlugin_logic_process_target_b = {{19{_zz_EU0_BranchPlugin_logic_process_target_b_2[12]}}, _zz_EU0_BranchPlugin_logic_process_target_b_2};
      end
    endcase
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
    EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE[0] = 1'b0;
  end

  assign EU0_BranchPlugin_logic_process_slices = (_zz_EU0_BranchPlugin_logic_process_slices + {1'b0,1'b1});
  assign EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE = (EU0_ExecutionUnitBase_pipeline_execute_0_PC + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_PC_TARGET = (EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND ? EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE : EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE);
  assign AguPlugin_logic_func3 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[14 : 12];
  assign when_AguPlugin_l89 = (EU0_ExecutionUnitBase_pipeline_execute_0_ready || EU0_ExecutionUnitBase_pipeline_execute_0_isRemoved);
  assign AguPlugin_setup_port_valid = ((EU0_ExecutionUnitBase_pipeline_execute_0_valid && EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SEL) && (! AguPlugin_logic_fired));
  assign AguPlugin_setup_port_payload_address = EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  assign AguPlugin_setup_port_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  assign AguPlugin_setup_port_payload_robIdMsb = EU0_ExecutionUnitBase_pipeline_execute_0_ROB_MSB;
  assign AguPlugin_setup_port_payload_size = AguPlugin_logic_func3[1 : 0];
  assign AguPlugin_setup_port_payload_sc = EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SC;
  assign AguPlugin_setup_port_payload_amo = EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_AMO;
  assign AguPlugin_setup_port_payload_swap = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[27];
  assign AguPlugin_setup_port_payload_op = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 29];
  assign AguPlugin_setup_port_payload_physicalRd = EU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  assign AguPlugin_setup_port_payload_writeRd = EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
  assign AguPlugin_setup_port_payload_aguId = EU0_ExecutionUnitBase_pipeline_execute_0_LSU_ID;
  assign AguPlugin_setup_port_payload_unsigned = AguPlugin_logic_func3[2];
  assign AguPlugin_setup_port_payload_pc = EU0_ExecutionUnitBase_pipeline_execute_0_PC;
  assign AguPlugin_setup_port_payload_lr = EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LR;
  assign AguPlugin_setup_port_payload_load = EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LOAD;
  assign AguPlugin_setup_port_payload_data = EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2;
  assign EU0_CsrAccessPlugin_setup_intFormatPort_valid = EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL;
  assign EU0_CsrAccessPlugin_logic_wake_wakeRobsSel = EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL;
  assign EU0_CsrAccessPlugin_logic_wake_wakeRegFileSel = EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL;
  always @(*) begin
    LsuPlugin_peripheralBus_cmd_ready = 1'b1;
    if(when_Stream_l1058) begin
      LsuPlugin_peripheralBus_cmd_ready = 1'b0;
    end
    if(when_Stream_l1058_1) begin
      LsuPlugin_peripheralBus_cmd_ready = 1'b0;
    end
  end

  assign when_Stream_l1058 = ((! LsuPlugin_peripheralBus_toAxiLite4_a_ready) && LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_0);
  assign when_Stream_l1058_1 = ((! LsuPlugin_peripheralBus_toAxiLite4_wRaw_ready) && LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_1);
  assign LsuPlugin_peripheralBus_toAxiLite4_a_valid = (LsuPlugin_peripheralBus_cmd_valid && LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_0);
  assign LsuPlugin_peripheralBus_toAxiLite4_a_payload_write = LsuPlugin_peripheralBus_cmd_payload_write;
  assign LsuPlugin_peripheralBus_toAxiLite4_a_payload_address = LsuPlugin_peripheralBus_cmd_payload_address;
  assign LsuPlugin_peripheralBus_toAxiLite4_a_payload_data = LsuPlugin_peripheralBus_cmd_payload_data;
  assign LsuPlugin_peripheralBus_toAxiLite4_a_payload_mask = LsuPlugin_peripheralBus_cmd_payload_mask;
  assign LsuPlugin_peripheralBus_toAxiLite4_a_payload_size = LsuPlugin_peripheralBus_cmd_payload_size;
  assign LsuPlugin_peripheralBus_toAxiLite4_a_fire = (LsuPlugin_peripheralBus_toAxiLite4_a_valid && LsuPlugin_peripheralBus_toAxiLite4_a_ready);
  assign LsuPlugin_peripheralBus_toAxiLite4_wRaw_valid = (LsuPlugin_peripheralBus_cmd_valid && LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_1);
  assign LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_write = LsuPlugin_peripheralBus_cmd_payload_write;
  assign LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_address = LsuPlugin_peripheralBus_cmd_payload_address;
  assign LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_data = LsuPlugin_peripheralBus_cmd_payload_data;
  assign LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_mask = LsuPlugin_peripheralBus_cmd_payload_mask;
  assign LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_size = LsuPlugin_peripheralBus_cmd_payload_size;
  assign LsuPlugin_peripheralBus_toAxiLite4_wRaw_fire = (LsuPlugin_peripheralBus_toAxiLite4_wRaw_valid && LsuPlugin_peripheralBus_toAxiLite4_wRaw_ready);
  assign when_Stream_l439 = (! LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_write);
  always @(*) begin
    LsuPlugin_peripheralBus_toAxiLite4_w_valid = LsuPlugin_peripheralBus_toAxiLite4_wRaw_valid;
    if(when_Stream_l439) begin
      LsuPlugin_peripheralBus_toAxiLite4_w_valid = 1'b0;
    end
  end

  always @(*) begin
    LsuPlugin_peripheralBus_toAxiLite4_wRaw_ready = LsuPlugin_peripheralBus_toAxiLite4_w_ready;
    if(when_Stream_l439) begin
      LsuPlugin_peripheralBus_toAxiLite4_wRaw_ready = 1'b1;
    end
  end

  assign LsuPlugin_peripheralBus_toAxiLite4_w_payload_write = LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_write;
  assign LsuPlugin_peripheralBus_toAxiLite4_w_payload_address = LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_address;
  assign LsuPlugin_peripheralBus_toAxiLite4_w_payload_data = LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_data;
  assign LsuPlugin_peripheralBus_toAxiLite4_w_payload_mask = LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_mask;
  assign LsuPlugin_peripheralBus_toAxiLite4_w_payload_size = LsuPlugin_peripheralBus_toAxiLite4_wRaw_payload_size;
  assign LsuPlugin_peripheralBus_toAxiLite4_a_ready = (LsuPlugin_peripheralBus_toAxiLite4_a_payload_write ? pBus_awready : pBus_arready);
  assign LsuPlugin_peripheralBus_toAxiLite4_addr = _zz_LsuPlugin_peripheralBus_toAxiLite4_addr;
  assign pBus_arvalid = (LsuPlugin_peripheralBus_toAxiLite4_a_valid && (! LsuPlugin_peripheralBus_toAxiLite4_a_payload_write));
  assign pBus_araddr = LsuPlugin_peripheralBus_toAxiLite4_addr;
  assign pBus_arprot = ((3'b000 | 3'b000) | 3'b000);
  assign pBus_awvalid = (LsuPlugin_peripheralBus_toAxiLite4_a_valid && LsuPlugin_peripheralBus_toAxiLite4_a_payload_write);
  assign pBus_awaddr = LsuPlugin_peripheralBus_toAxiLite4_addr;
  assign pBus_awprot = ((3'b000 | 3'b000) | 3'b000);
  assign pBus_wvalid = LsuPlugin_peripheralBus_toAxiLite4_w_valid;
  assign pBus_wdata = LsuPlugin_peripheralBus_toAxiLite4_w_payload_data;
  assign pBus_wstrb = LsuPlugin_peripheralBus_toAxiLite4_w_payload_mask;
  assign LsuPlugin_peripheralBus_toAxiLite4_w_ready = pBus_wready;
  assign LsuPlugin_peripheralBus_rsp_valid = (pBus_rvalid || pBus_bvalid);
  assign LsuPlugin_peripheralBus_rsp_payload_data = pBus_rdata;
  assign LsuPlugin_peripheralBus_rsp_payload_error = (! (LsuPlugin_peripheralBus_toAxiLite4_writeSel ? (pBus_bresp == 2'b00) : (pBus_rresp == 2'b00)));
  assign pBus_bready = 1'b1;
  assign pBus_rready = 1'b1;
  assign dBusAxi_arvalid = DataCachePlugin_mem_read_cmd_valid;
  assign dBusAxi_araddr = DataCachePlugin_mem_read_cmd_payload_address;
  assign dBusAxi_arid = DataCachePlugin_mem_read_cmd_payload_id;
  assign dBusAxi_arprot = 3'b010;
  assign dBusAxi_arlen = 8'h0f;
  assign dBusAxi_arsize = 3'b010;
  assign dBusAxi_arburst = 2'b01;
  assign DataCachePlugin_mem_read_cmd_ready = dBusAxi_arready;
  assign DataCachePlugin_mem_read_rsp_valid = dBusAxi_rvalid;
  assign DataCachePlugin_mem_read_rsp_payload_data = dBusAxi_rdata;
  assign DataCachePlugin_mem_read_rsp_payload_id = dBusAxi_rid;
  assign DataCachePlugin_mem_read_rsp_payload_error = (! (dBusAxi_rresp == 2'b00));
  assign dBusAxi_rready = 1'b1;
  always @(*) begin
    DataCachePlugin_mem_write_cmd_ready = 1'b1;
    if(when_Stream_l1058_2) begin
      DataCachePlugin_mem_write_cmd_ready = 1'b0;
    end
    if(when_Stream_l1058_3) begin
      DataCachePlugin_mem_write_cmd_ready = 1'b0;
    end
  end

  assign when_Stream_l1058_2 = ((! DataCachePlugin_mem_toAxi4_awRaw_ready) && DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_0);
  assign when_Stream_l1058_3 = ((! DataCachePlugin_mem_toAxi4_wRaw_ready) && DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_1);
  assign DataCachePlugin_mem_toAxi4_awRaw_valid = (DataCachePlugin_mem_write_cmd_valid && DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_0);
  assign DataCachePlugin_mem_toAxi4_awRaw_payload_last = DataCachePlugin_mem_write_cmd_payload_last;
  assign DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_address = DataCachePlugin_mem_write_cmd_payload_fragment_address;
  assign DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_data = DataCachePlugin_mem_write_cmd_payload_fragment_data;
  assign DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_id = DataCachePlugin_mem_write_cmd_payload_fragment_id;
  assign DataCachePlugin_mem_toAxi4_awRaw_fire = (DataCachePlugin_mem_toAxi4_awRaw_valid && DataCachePlugin_mem_toAxi4_awRaw_ready);
  assign DataCachePlugin_mem_toAxi4_wRaw_valid = (DataCachePlugin_mem_write_cmd_valid && DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_1);
  assign DataCachePlugin_mem_toAxi4_wRaw_payload_last = DataCachePlugin_mem_write_cmd_payload_last;
  assign DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_address = DataCachePlugin_mem_write_cmd_payload_fragment_address;
  assign DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_data = DataCachePlugin_mem_write_cmd_payload_fragment_data;
  assign DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_id = DataCachePlugin_mem_write_cmd_payload_fragment_id;
  assign DataCachePlugin_mem_toAxi4_wRaw_fire = (DataCachePlugin_mem_toAxi4_wRaw_valid && DataCachePlugin_mem_toAxi4_wRaw_ready);
  assign when_Stream_l439_1 = (! DataCachePlugin_mem_toAxi4_awRaw_payload_first);
  always @(*) begin
    DataCachePlugin_mem_toAxi4_awFiltred_valid = DataCachePlugin_mem_toAxi4_awRaw_valid;
    if(when_Stream_l439_1) begin
      DataCachePlugin_mem_toAxi4_awFiltred_valid = 1'b0;
    end
  end

  always @(*) begin
    DataCachePlugin_mem_toAxi4_awRaw_ready = DataCachePlugin_mem_toAxi4_awFiltred_ready;
    if(when_Stream_l439_1) begin
      DataCachePlugin_mem_toAxi4_awRaw_ready = 1'b1;
    end
  end

  assign DataCachePlugin_mem_toAxi4_awFiltred_payload_last = DataCachePlugin_mem_toAxi4_awRaw_payload_last;
  assign DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_address = DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_address;
  assign DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_data = DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_data;
  assign DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_id = DataCachePlugin_mem_toAxi4_awRaw_payload_fragment_id;
  always @(*) begin
    DataCachePlugin_mem_toAxi4_awFiltred_ready = DataCachePlugin_mem_toAxi4_aw_ready;
    if(when_Stream_l369_1) begin
      DataCachePlugin_mem_toAxi4_awFiltred_ready = 1'b1;
    end
  end

  assign when_Stream_l369_1 = (! DataCachePlugin_mem_toAxi4_aw_valid);
  assign DataCachePlugin_mem_toAxi4_aw_valid = DataCachePlugin_mem_toAxi4_awFiltred_rValid;
  assign DataCachePlugin_mem_toAxi4_aw_payload_last = DataCachePlugin_mem_toAxi4_awFiltred_rData_last;
  assign DataCachePlugin_mem_toAxi4_aw_payload_fragment_address = DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_address;
  assign DataCachePlugin_mem_toAxi4_aw_payload_fragment_data = DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_data;
  assign DataCachePlugin_mem_toAxi4_aw_payload_fragment_id = DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_id;
  assign dBusAxi_awvalid = DataCachePlugin_mem_toAxi4_aw_valid;
  assign dBusAxi_awaddr = DataCachePlugin_mem_toAxi4_aw_payload_fragment_address;
  assign dBusAxi_awid = DataCachePlugin_mem_toAxi4_aw_payload_fragment_id;
  assign dBusAxi_awprot = 3'b010;
  assign dBusAxi_awlen = 8'h0f;
  assign dBusAxi_awsize = 3'b010;
  assign dBusAxi_awburst = 2'b01;
  assign DataCachePlugin_mem_toAxi4_aw_ready = dBusAxi_awready;
  assign _zz_DataCachePlugin_mem_toAxi4_wRaw_ready = (! DataCachePlugin_mem_toAxi4_awFiltred_valid);
  assign DataCachePlugin_mem_toAxi4_w_valid = (DataCachePlugin_mem_toAxi4_wRaw_valid && _zz_DataCachePlugin_mem_toAxi4_wRaw_ready);
  assign DataCachePlugin_mem_toAxi4_wRaw_ready = (DataCachePlugin_mem_toAxi4_w_ready && _zz_DataCachePlugin_mem_toAxi4_wRaw_ready);
  assign DataCachePlugin_mem_toAxi4_w_payload_last = DataCachePlugin_mem_toAxi4_wRaw_payload_last;
  assign DataCachePlugin_mem_toAxi4_w_payload_fragment_address = DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_address;
  assign DataCachePlugin_mem_toAxi4_w_payload_fragment_data = DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_data;
  assign DataCachePlugin_mem_toAxi4_w_payload_fragment_id = DataCachePlugin_mem_toAxi4_wRaw_payload_fragment_id;
  assign dBusAxi_wvalid = DataCachePlugin_mem_toAxi4_w_valid;
  assign dBusAxi_wdata = DataCachePlugin_mem_toAxi4_w_payload_fragment_data;
  assign dBusAxi_wstrb = 4'b1111;
  assign dBusAxi_wlast = DataCachePlugin_mem_toAxi4_w_payload_last;
  assign DataCachePlugin_mem_toAxi4_w_ready = dBusAxi_wready;
  assign DataCachePlugin_mem_write_rsp_valid = dBusAxi_bvalid;
  assign DataCachePlugin_mem_write_rsp_payload_id = dBusAxi_bid;
  assign DataCachePlugin_mem_write_rsp_payload_error = (! (dBusAxi_bresp == 2'b00));
  assign dBusAxi_bready = 1'b1;
  assign PrivilegedPlugin_io_int_machine_external = plicCtrl_io_targets[0];
  assign PrivilegedPlugin_io_int_machine_timer = clintCtrl_io_timerInterrupt[0];
  assign PrivilegedPlugin_io_int_machine_software = clintCtrl_io_softwareInterrupt[0];
  assign PrivilegedPlugin_io_int_supervisor_external = plicCtrl_io_targets[1];
  assign PrivilegedPlugin_io_rdtime = clintCtrl_io_time;
  assign FrontendPlugin_allocated_haltRequest_FrontendPlugin_l67 = CommitPlugin_logic_reschedule_valid;
  always @(*) begin
    integer_RfTranslationPlugin_logic_impl_io_rollback = CommitPlugin_logic_commit_reschedulePort_valid;
    if(integer_RfTranslationPlugin_logic_init_busy) begin
      integer_RfTranslationPlugin_logic_impl_io_rollback = 1'b1;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_writes_0_valid = (((FrontendPlugin_allocated_isFireing && FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0) && FrontendPlugin_allocated_WRITE_RD_0) && 1'b1);
  always @(*) begin
    integer_RfTranslationPlugin_logic_impl_io_commits_0_valid = ((CommitPlugin_logic_commit_event_mask[0] && integer_RfTranslationPlugin_logic_onCommit_writeRd_0) && 1'b1);
    if(integer_RfTranslationPlugin_logic_init_busy) begin
      integer_RfTranslationPlugin_logic_impl_io_commits_0_valid = 1'b1;
    end
  end

  always @(*) begin
    integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_address = integer_RfTranslationPlugin_logic_onCommit_archRd_0;
    if(integer_RfTranslationPlugin_logic_init_busy) begin
      integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_address = integer_RfTranslationPlugin_logic_init_counter[4:0];
    end
  end

  always @(*) begin
    integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_data = integer_RfTranslationPlugin_logic_onCommit_physRd_0;
    if(integer_RfTranslationPlugin_logic_init_busy) begin
      integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_data = 6'h00;
    end
  end

  assign integer_RfTranslationPlugin_logic_init_busy = (! integer_RfTranslationPlugin_logic_init_counter[5]);
  assign when_RfTranslationPlugin_l193 = 1'b1;
  assign integer_RfTranslationPlugin_logic_impl_io_reads_0_cmd_valid = (FrontendPlugin_allocated_WRITE_RD_0 && when_RfTranslationPlugin_l193);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RD_FREE_0 = 6'bxxxxxx;
    if(when_RfTranslationPlugin_l193) begin
      FrontendPlugin_allocated_PHYS_RD_FREE_0 = integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_payload;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_reads_1_cmd_valid = (FrontendPlugin_allocated_READ_RS_0_0 && 1'b1);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RS_0_0 = 6'bxxxxxx;
    if(1'b1) begin
      FrontendPlugin_allocated_PHYS_RS_0_0 = integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_payload;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_reads_2_cmd_valid = (FrontendPlugin_allocated_READ_RS_1_0 && 1'b1);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RS_1_0 = 6'bxxxxxx;
    if(1'b1) begin
      FrontendPlugin_allocated_PHYS_RS_1_0 = integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_payload;
    end
  end

  always @(*) begin
    integer_RfAllocationPlugin_logic_allocator_io_push_0_valid = (((CommitPlugin_logic_free_port_valid && integer_RfAllocationPlugin_logic_push_mask_0) && integer_RfAllocationPlugin_logic_push_writeRd_0) && 1'b1);
    if(when_RfAllocationPlugin_l81) begin
      integer_RfAllocationPlugin_logic_allocator_io_push_0_valid = 1'b0;
    end
    if(integer_RfAllocationPlugin_logic_init_busy) begin
      integer_RfAllocationPlugin_logic_allocator_io_push_0_valid = 1'b1;
    end
  end

  always @(*) begin
    integer_RfAllocationPlugin_logic_allocator_io_push_0_payload = (CommitPlugin_logic_free_port_payload_commited[0] ? integer_RfAllocationPlugin_logic_push_physicalRdOld_0 : integer_RfAllocationPlugin_logic_push_physicalRdNew_0);
    if(integer_RfAllocationPlugin_logic_init_busy) begin
      integer_RfAllocationPlugin_logic_allocator_io_push_0_payload = integer_RfAllocationPlugin_logic_init_counter[5:0];
    end
  end

  assign when_RfAllocationPlugin_l81 = (integer_RfAllocationPlugin_logic_allocator_io_push_0_payload == 6'h00);
  assign integer_RfAllocationPlugin_logic_init_busy = (! integer_RfAllocationPlugin_logic_init_counter[6]);
  assign BranchContextPlugin_logic_onCommit_isBranchCommit_0 = (CommitPlugin_logic_commit_event_mask[0] && BranchContextPlugin_logic_onCommit_isBranch_0);
  assign BranchContextPlugin_logic_onCommit_commitedNext = (BranchContextPlugin_logic_ptr_commited + _zz_BranchContextPlugin_logic_onCommit_commitedNext);
  assign HistoryPlugin_logic_onCommit_valueNext = HistoryPlugin_logic_onCommit_value;
  assign HistoryPlugin_logic_onCommit_whitebox_0 = HistoryPlugin_logic_onCommit_valueNext;
  assign when_HistoryPlugin_l90 = (CommitPlugin_logic_commit_event_mask[0] && HistoryPlugin_logic_onCommit_isConditionalBranch_0);
  always @(*) begin
    HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_value;
    if(BtbPlugin_setup_historyPush_flush) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_update_pushes_0_stateNext_1;
    end
    if(FetchCachePlugin_setup_historyJump_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = FetchCachePlugin_setup_historyJump_payload_history;
    end
    if(DecoderPredictionPlugin_setup_historyPush_flush) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_update_pushes_2_stateNext_1;
    end
    if(CommitPlugin_logic_reschedule_reschedulePort_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_update_rescheduleFlush_newHistory;
    end
  end

  assign FetchPlugin_stages_0_BRANCH_HISTORY = HistoryPlugin_logic_onFetch_valueNext;
  assign HistoryPlugin_logic_update_pushes_0_stateNext = HistoryPlugin_logic_update_pushes_0_state;
  assign when_HistoryPlugin_l115 = BtbPlugin_setup_historyPush_mask[0];
  assign HistoryPlugin_logic_update_pushes_2_stateNext = HistoryPlugin_logic_update_pushes_2_state;
  assign when_HistoryPlugin_l115_1 = DecoderPredictionPlugin_setup_historyPush_mask[0];
  assign HistoryPlugin_logic_update_rescheduleFlush_instHistory = _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_1[23 : 0];
  assign HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch = _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_1[0];
  assign HistoryPlugin_logic_update_rescheduleFlush_isTaken = _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_1[0];
  assign HistoryPlugin_logic_update_rescheduleFlush_newHistory = (HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch ? {HistoryPlugin_logic_update_rescheduleFlush_instHistory[22 : 0],HistoryPlugin_logic_update_rescheduleFlush_isTaken} : HistoryPlugin_logic_update_rescheduleFlush_instHistory);
  assign DecoderPredictionPlugin_logic_ras_healPush = _zz_DecoderPredictionPlugin_logic_ras_healPush_1[3 : 0];
  assign DecoderPredictionPlugin_logic_ras_healPop = (DecoderPredictionPlugin_logic_ras_healPush - 4'b0001);
  assign DecoderPredictionPlugin_logic_decodePatch_rasPushUsed = 1'b0;
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          3'b000 : begin
            Lsu2Plugin_logic_lq_regs_0_allocation = 1'b1;
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315) begin
      Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_2)
          3'b000 : begin
            Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b1;
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_118) begin
          Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_118) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_delete = 1'b0;
    if(when_Lsu2Plugin_l454) begin
      Lsu2Plugin_logic_lq_regs_0_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_0_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_118) begin
            Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_118) begin
              Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_118) begin
            Lsu2Plugin_logic_lq_regs_0_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_118) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315 = ((((|(Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_0_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_0_waitOn_sqId)));
  assign when_Lsu2Plugin_l338 = (Lsu2Plugin_logic_lq_regs_0_redoSet || Lsu2Plugin_logic_lq_regs_0_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
            Lsu2Plugin_logic_lq_regs_1_allocation = 1'b1;
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_1) begin
      Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_2)
          3'b000 : begin
          end
          3'b001 : begin
            Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b1;
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_119) begin
          Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_119) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_delete = 1'b0;
    if(when_Lsu2Plugin_l454_1) begin
      Lsu2Plugin_logic_lq_regs_1_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_1_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_119) begin
            Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_119) begin
              Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_119) begin
            Lsu2Plugin_logic_lq_regs_1_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_119) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_1 = ((((|(Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_1_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_1_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_1 = (Lsu2Plugin_logic_lq_regs_1_redoSet || Lsu2Plugin_logic_lq_regs_1_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
            Lsu2Plugin_logic_lq_regs_2_allocation = 1'b1;
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_2) begin
      Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_2)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
            Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b1;
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_120) begin
          Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_120) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_delete = 1'b0;
    if(when_Lsu2Plugin_l454_2) begin
      Lsu2Plugin_logic_lq_regs_2_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_2_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_120) begin
            Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_120) begin
              Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_120) begin
            Lsu2Plugin_logic_lq_regs_2_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_120) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_2 = ((((|(Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_2_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_2_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_2 = (Lsu2Plugin_logic_lq_regs_2_redoSet || Lsu2Plugin_logic_lq_regs_2_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
            Lsu2Plugin_logic_lq_regs_3_allocation = 1'b1;
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_3) begin
      Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_2)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
            Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b1;
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_121) begin
          Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_121) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_delete = 1'b0;
    if(when_Lsu2Plugin_l454_3) begin
      Lsu2Plugin_logic_lq_regs_3_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_3_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_121) begin
            Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_121) begin
              Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_121) begin
            Lsu2Plugin_logic_lq_regs_3_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_121) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_3 = ((((|(Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_3_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_3_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_3 = (Lsu2Plugin_logic_lq_regs_3_redoSet || Lsu2Plugin_logic_lq_regs_3_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
            Lsu2Plugin_logic_lq_regs_4_allocation = 1'b1;
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_4) begin
      Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_2)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
            Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b1;
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_122) begin
          Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_122) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_delete = 1'b0;
    if(when_Lsu2Plugin_l454_4) begin
      Lsu2Plugin_logic_lq_regs_4_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_4_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_122) begin
            Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_122) begin
              Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_122) begin
            Lsu2Plugin_logic_lq_regs_4_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_122) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_4 = ((((|(Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_4_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_4_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_4 = (Lsu2Plugin_logic_lq_regs_4_redoSet || Lsu2Plugin_logic_lq_regs_4_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
            Lsu2Plugin_logic_lq_regs_5_allocation = 1'b1;
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_5) begin
      Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_2)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
            Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b1;
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_123) begin
          Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_123) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_delete = 1'b0;
    if(when_Lsu2Plugin_l454_5) begin
      Lsu2Plugin_logic_lq_regs_5_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_5_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_123) begin
            Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_123) begin
              Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_123) begin
            Lsu2Plugin_logic_lq_regs_5_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_123) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_5 = ((((|(Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_5_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_5_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_5 = (Lsu2Plugin_logic_lq_regs_5_redoSet || Lsu2Plugin_logic_lq_regs_5_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
            Lsu2Plugin_logic_lq_regs_6_allocation = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_6) begin
      Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_2)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
            Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_124) begin
          Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_124) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_delete = 1'b0;
    if(when_Lsu2Plugin_l454_6) begin
      Lsu2Plugin_logic_lq_regs_6_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_6_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_124) begin
            Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_124) begin
              Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_124) begin
            Lsu2Plugin_logic_lq_regs_6_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_124) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_6 = ((((|(Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_6_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_6_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_6 = (Lsu2Plugin_logic_lq_regs_6_redoSet || Lsu2Plugin_logic_lq_regs_6_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
            Lsu2Plugin_logic_lq_regs_7_allocation = 1'b1;
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_7) begin
      Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_2)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
            Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b1;
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_125) begin
          Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_125) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_delete = 1'b0;
    if(when_Lsu2Plugin_l454_7) begin
      Lsu2Plugin_logic_lq_regs_7_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_7_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_125) begin
            Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_125) begin
              Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_125) begin
            Lsu2Plugin_logic_lq_regs_7_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_125) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_7 = ((((|(Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_7_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_7_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_7 = (Lsu2Plugin_logic_lq_regs_7_redoSet || Lsu2Plugin_logic_lq_regs_7_delete);
  assign Lsu2Plugin_logic_lq_ptr_allocReal = Lsu2Plugin_logic_lq_ptr_alloc[2 : 0];
  assign Lsu2Plugin_logic_lq_ptr_freeReal = Lsu2Plugin_logic_lq_ptr_free[2 : 0];
  assign when_UInt_l120 = (|Lsu2Plugin_logic_lq_tracker_freeNext[3 : 1]);
  always @(*) begin
    if(when_UInt_l120) begin
      _zz_Lsu2Plugin_logic_lq_tracker_freeReduced = 1'b1;
    end else begin
      _zz_Lsu2Plugin_logic_lq_tracker_freeReduced = Lsu2Plugin_logic_lq_tracker_freeNext[0 : 0];
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_tracker_freeNext = (_zz_Lsu2Plugin_logic_lq_tracker_freeNext - _zz_Lsu2Plugin_logic_lq_tracker_freeNext_2);
    if(Lsu2Plugin_logic_lq_tracker_clear) begin
      Lsu2Plugin_logic_lq_tracker_freeNext = 4'b1000;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_tracker_clear = 1'b0;
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_tracker_clear = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_lq_onCommit_lqCommits_0 = (CommitPlugin_logic_commit_event_mask[0] && Lsu2Plugin_logic_lq_onCommit_lqAlloc_0);
  assign Lsu2Plugin_logic_lq_onCommit_lqCommitCount = _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount;
  assign Lsu2Plugin_logic_lq_onCommit_free = Lsu2Plugin_logic_lq_ptr_free;
  assign Lsu2Plugin_logic_lq_onCommit_priority = Lsu2Plugin_logic_lq_ptr_priority;
  assign when_Lsu2Plugin_l454 = ((_zz_when_Lsu2Plugin_l454 == 3'b000) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_1 = ((_zz_when_Lsu2Plugin_l454_1 == 3'b001) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_2 = ((_zz_when_Lsu2Plugin_l454_2 == 3'b010) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_3 = ((_zz_when_Lsu2Plugin_l454_3 == 3'b011) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_4 = ((_zz_when_Lsu2Plugin_l454_4 == 3'b100) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_5 = ((_zz_when_Lsu2Plugin_l454_5 == 3'b101) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_6 = ((_zz_when_Lsu2Plugin_l454_6 == 3'b110) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_7 = ((_zz_when_Lsu2Plugin_l454_7 == 3'b111) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign Lsu2Plugin_logic_lq_tracker_add = Lsu2Plugin_logic_lq_onCommit_lqCommitCount;
  always @(*) begin
    Lsu2Plugin_logic_lq_reservation_kill = 1'b0;
    if(DataCachePlugin_setup_writebackBusy) begin
      Lsu2Plugin_logic_lq_reservation_kill = 1'b1;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
        if(when_Lsu2Plugin_l1715) begin
          Lsu2Plugin_logic_lq_reservation_kill = 1'b1;
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign when_Lsu2Plugin_l484 = Lsu2Plugin_logic_lq_reservation_counter[6];
  assign Lsu2Plugin_logic_lq_hazardPrediction_hazard = 1'b0;
  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_valid = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_VALID;
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_valid = 1'b1;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address = 7'bxxxxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC[8 : 2];
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC[8 : 2];
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'bxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE + _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score);
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'b111;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag = 16'bxxxxxxxxxxxxxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC[24 : 9];
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC[24 : 9];
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta = 3'bxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_DELTA;
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta = _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta[2:0];
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_valid = (Lsu2Plugin_logic_lq_hazardPrediction_write_valid && (! Lsu2Plugin_logic_lq_hazardPrediction_hazard));
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_address = Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address;
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_score = Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score;
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_tag = Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag;
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_delta = Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta;
  assign Lsu2Plugin_logic_lq_hitPrediction_hazard = 1'b0;
  assign Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_valid = (Lsu2Plugin_logic_lq_hitPrediction_write_valid && (! Lsu2Plugin_logic_lq_hitPrediction_hazard));
  assign Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_address = Lsu2Plugin_logic_lq_hitPrediction_write_payload_address;
  assign Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_data_counter = Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter;
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          3'b000 : begin
            Lsu2Plugin_logic_sq_regs_0_allocation = 1'b1;
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369) begin
      Lsu2Plugin_logic_sq_regs_0_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_3)
          3'b000 : begin
            Lsu2Plugin_logic_sq_regs_0_redoSet = 1'b1;
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_126) begin
          Lsu2Plugin_logic_sq_regs_0_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524) begin
        Lsu2Plugin_logic_sq_regs_0_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1913) begin
        Lsu2Plugin_logic_sq_regs_0_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_commitedNext = Lsu2Plugin_logic_sq_regs_0_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_44[0]) begin
        Lsu2Plugin_logic_sq_regs_0_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_126) begin
              Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369 = (Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385 = (Lsu2Plugin_logic_sq_regs_0_redoSet || Lsu2Plugin_logic_sq_regs_0_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
            Lsu2Plugin_logic_sq_regs_1_allocation = 1'b1;
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_1) begin
      Lsu2Plugin_logic_sq_regs_1_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_3)
          3'b000 : begin
          end
          3'b001 : begin
            Lsu2Plugin_logic_sq_regs_1_redoSet = 1'b1;
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_127) begin
          Lsu2Plugin_logic_sq_regs_1_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_1) begin
        Lsu2Plugin_logic_sq_regs_1_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1913_1) begin
        Lsu2Plugin_logic_sq_regs_1_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_commitedNext = Lsu2Plugin_logic_sq_regs_1_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_44[1]) begin
        Lsu2Plugin_logic_sq_regs_1_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_127) begin
              Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_1 = (Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_1 = (Lsu2Plugin_logic_sq_regs_1_redoSet || Lsu2Plugin_logic_sq_regs_1_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
            Lsu2Plugin_logic_sq_regs_2_allocation = 1'b1;
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_2) begin
      Lsu2Plugin_logic_sq_regs_2_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_3)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
            Lsu2Plugin_logic_sq_regs_2_redoSet = 1'b1;
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_128) begin
          Lsu2Plugin_logic_sq_regs_2_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_2) begin
        Lsu2Plugin_logic_sq_regs_2_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1913_2) begin
        Lsu2Plugin_logic_sq_regs_2_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_commitedNext = Lsu2Plugin_logic_sq_regs_2_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_44[2]) begin
        Lsu2Plugin_logic_sq_regs_2_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_128) begin
              Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_2 = (Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_2 = (Lsu2Plugin_logic_sq_regs_2_redoSet || Lsu2Plugin_logic_sq_regs_2_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
            Lsu2Plugin_logic_sq_regs_3_allocation = 1'b1;
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_3) begin
      Lsu2Plugin_logic_sq_regs_3_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_3)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
            Lsu2Plugin_logic_sq_regs_3_redoSet = 1'b1;
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_129) begin
          Lsu2Plugin_logic_sq_regs_3_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_3) begin
        Lsu2Plugin_logic_sq_regs_3_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1913_3) begin
        Lsu2Plugin_logic_sq_regs_3_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_commitedNext = Lsu2Plugin_logic_sq_regs_3_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_44[3]) begin
        Lsu2Plugin_logic_sq_regs_3_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_129) begin
              Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_3 = (Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_3 = (Lsu2Plugin_logic_sq_regs_3_redoSet || Lsu2Plugin_logic_sq_regs_3_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
            Lsu2Plugin_logic_sq_regs_4_allocation = 1'b1;
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_4) begin
      Lsu2Plugin_logic_sq_regs_4_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_3)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
            Lsu2Plugin_logic_sq_regs_4_redoSet = 1'b1;
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_130) begin
          Lsu2Plugin_logic_sq_regs_4_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_4) begin
        Lsu2Plugin_logic_sq_regs_4_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1913_4) begin
        Lsu2Plugin_logic_sq_regs_4_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_commitedNext = Lsu2Plugin_logic_sq_regs_4_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_44[4]) begin
        Lsu2Plugin_logic_sq_regs_4_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_130) begin
              Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_4 = (Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_4 = (Lsu2Plugin_logic_sq_regs_4_redoSet || Lsu2Plugin_logic_sq_regs_4_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
            Lsu2Plugin_logic_sq_regs_5_allocation = 1'b1;
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_5) begin
      Lsu2Plugin_logic_sq_regs_5_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_3)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
            Lsu2Plugin_logic_sq_regs_5_redoSet = 1'b1;
          end
          3'b110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_131) begin
          Lsu2Plugin_logic_sq_regs_5_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_5) begin
        Lsu2Plugin_logic_sq_regs_5_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1913_5) begin
        Lsu2Plugin_logic_sq_regs_5_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_commitedNext = Lsu2Plugin_logic_sq_regs_5_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_44[5]) begin
        Lsu2Plugin_logic_sq_regs_5_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_131) begin
              Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_5 = (Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_5 = (Lsu2Plugin_logic_sq_regs_5_redoSet || Lsu2Plugin_logic_sq_regs_5_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
            Lsu2Plugin_logic_sq_regs_6_allocation = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_6) begin
      Lsu2Plugin_logic_sq_regs_6_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_3)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
            Lsu2Plugin_logic_sq_regs_6_redoSet = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_132) begin
          Lsu2Plugin_logic_sq_regs_6_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_6) begin
        Lsu2Plugin_logic_sq_regs_6_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1913_6) begin
        Lsu2Plugin_logic_sq_regs_6_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_commitedNext = Lsu2Plugin_logic_sq_regs_6_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_44[6]) begin
        Lsu2Plugin_logic_sq_regs_6_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_132) begin
              Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_6 = (Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_6 = (Lsu2Plugin_logic_sq_regs_6_redoSet || Lsu2Plugin_logic_sq_regs_6_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
            Lsu2Plugin_logic_sq_regs_7_allocation = 1'b1;
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_7) begin
      Lsu2Plugin_logic_sq_regs_7_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1423_3)
          3'b000 : begin
          end
          3'b001 : begin
          end
          3'b010 : begin
          end
          3'b011 : begin
          end
          3'b100 : begin
          end
          3'b101 : begin
          end
          3'b110 : begin
          end
          default : begin
            Lsu2Plugin_logic_sq_regs_7_redoSet = 1'b1;
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_133) begin
          Lsu2Plugin_logic_sq_regs_7_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_7) begin
        Lsu2Plugin_logic_sq_regs_7_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1913_7) begin
        Lsu2Plugin_logic_sq_regs_7_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_commitedNext = Lsu2Plugin_logic_sq_regs_7_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_44[7]) begin
        Lsu2Plugin_logic_sq_regs_7_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_133) begin
              Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_7 = (Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_7 = (Lsu2Plugin_logic_sq_regs_7_redoSet || Lsu2Plugin_logic_sq_regs_7_delete);
  assign Lsu2Plugin_logic_sq_ptr_allocReal = Lsu2Plugin_logic_sq_ptr_alloc[2 : 0];
  assign Lsu2Plugin_logic_sq_ptr_freeReal = Lsu2Plugin_logic_sq_ptr_free[2 : 0];
  assign Lsu2Plugin_logic_sq_ptr_writeBackReal = Lsu2Plugin_logic_sq_ptr_writeBack[2 : 0];
  assign Lsu2Plugin_logic_sq_ptr_commitReal = Lsu2Plugin_logic_sq_ptr_commit[2 : 0];
  assign Lsu2Plugin_logic_sqWritebackEvent_valid = Lsu2Plugin_logic_sq_ptr_onFree_valid;
  assign Lsu2Plugin_logic_sqWritebackEvent_payload = Lsu2Plugin_logic_sq_ptr_onFree_payload;
  assign when_Lsu2Plugin_l572 = (Lsu2Plugin_logic_sq_ptr_commit != Lsu2Plugin_logic_sq_ptr_free);
  assign when_UInt_l120_1 = (|Lsu2Plugin_logic_sq_tracker_freeNext[3 : 1]);
  always @(*) begin
    if(when_UInt_l120_1) begin
      _zz_Lsu2Plugin_logic_sq_tracker_freeReduced = 1'b1;
    end else begin
      _zz_Lsu2Plugin_logic_sq_tracker_freeReduced = Lsu2Plugin_logic_sq_tracker_freeNext[0 : 0];
    end
  end

  assign Lsu2Plugin_logic_sq_tracker_freeNext = (_zz_Lsu2Plugin_logic_sq_tracker_freeNext + _zz_Lsu2Plugin_logic_sq_tracker_freeNext_4);
  assign Lsu2Plugin_logic_sq_onCommit_sqCommits_0 = (CommitPlugin_logic_commit_event_mask[0] && Lsu2Plugin_logic_sq_onCommit_sqAlloc_0);
  assign Lsu2Plugin_logic_sq_onCommit_commitComb = Lsu2Plugin_logic_sq_ptr_commit;
  assign when_Lsu2Plugin_l591 = (CommitPlugin_logic_commit_event_mask[0] && Lsu2Plugin_logic_sq_onCommit_sqAlloc_0);
  assign _zz_44 = ({7'd0,1'b1} <<< Lsu2Plugin_logic_sq_onCommit_commitComb[2 : 0]);
  assign Lsu2Plugin_logic_sq_ptr_commitNext = Lsu2Plugin_logic_sq_onCommit_commitComb_1;
  always @(*) begin
    FrontendPlugin_dispatch_LSU_ID_0 = 4'bxxxx;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      FrontendPlugin_dispatch_LSU_ID_0 = Lsu2Plugin_logic_allocation_loads_alloc;
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      FrontendPlugin_dispatch_LSU_ID_0 = Lsu2Plugin_logic_allocation_stores_alloc;
    end
  end

  assign Lsu2Plugin_logic_allocation_loads_requests_0 = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 && FrontendPlugin_dispatch_LQ_ALLOC_0);
  assign Lsu2Plugin_logic_allocation_loads_requestsCount = _zz_Lsu2Plugin_logic_allocation_loads_requestsCount;
  assign Lsu2Plugin_logic_allocation_loads_full = (Lsu2Plugin_logic_lq_tracker_freeReduced < Lsu2Plugin_logic_allocation_loads_requestsCount);
  assign Lsu2Plugin_logic_allocation_loads_alloc = Lsu2Plugin_logic_lq_ptr_alloc;
  assign Lsu2Plugin_logic_allocation_stores_requests_0 = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 && FrontendPlugin_dispatch_SQ_ALLOC_0);
  assign Lsu2Plugin_logic_allocation_stores_requestsCount = _zz_Lsu2Plugin_logic_allocation_stores_requestsCount;
  assign Lsu2Plugin_logic_allocation_stores_full = (Lsu2Plugin_logic_sq_tracker_freeReduced < Lsu2Plugin_logic_allocation_stores_requestsCount);
  assign Lsu2Plugin_logic_allocation_stores_alloc = Lsu2Plugin_logic_sq_ptr_alloc;
  assign FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l620 = (FrontendPlugin_dispatch_valid && (Lsu2Plugin_logic_allocation_loads_full || Lsu2Plugin_logic_allocation_stores_full));
  assign FrontendPlugin_dispatch_LQ_ID_0 = Lsu2Plugin_logic_allocation_loads_alloc[2:0];
  assign FrontendPlugin_dispatch_SQ_ID_0 = Lsu2Plugin_logic_allocation_stores_alloc[2:0];
  assign FrontendPlugin_dispatch_isFireing = (FrontendPlugin_dispatch_valid && FrontendPlugin_dispatch_ready);
  always @(*) begin
    Lsu2Plugin_logic_lq_tracker_sub = 1'b0;
    if(FrontendPlugin_dispatch_isFireing) begin
      Lsu2Plugin_logic_lq_tracker_sub = Lsu2Plugin_logic_allocation_loads_requestsCount;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_tracker_sub = 1'b0;
    if(FrontendPlugin_dispatch_isFireing) begin
      Lsu2Plugin_logic_sq_tracker_sub = Lsu2Plugin_logic_allocation_stores_requestsCount;
    end
  end

  assign Lsu2Plugin_logic_aguPush_0_pushLq = (AguPlugin_setup_port_valid && AguPlugin_setup_port_payload_load);
  assign Lsu2Plugin_logic_aguPush_0_pushSq = (AguPlugin_setup_port_valid && (! AguPlugin_setup_port_payload_load));
  always @(*) begin
    _zz_Lsu2Plugin_logic_aguPush_0_dataMask = 4'bxxxx;
    case(AguPlugin_setup_port_payload_size)
      2'b00 : begin
        _zz_Lsu2Plugin_logic_aguPush_0_dataMask = 4'b0001;
      end
      2'b01 : begin
        _zz_Lsu2Plugin_logic_aguPush_0_dataMask = 4'b0011;
      end
      2'b10 : begin
        _zz_Lsu2Plugin_logic_aguPush_0_dataMask = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_aguPush_0_dataMask = (_zz_Lsu2Plugin_logic_aguPush_0_dataMask <<< AguPlugin_setup_port_payload_address[1 : 0]);
  assign switch_Utils_l1423 = AguPlugin_setup_port_payload_aguId[2:0];
  assign _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score = Lsu2Plugin_logic_lq_hazardPrediction_mem_spinal_port1;
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score = _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score[2 : 0];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_tag = _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score[18 : 3];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_delta = _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score[21 : 19];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_valid = AguPlugin_setup_port_payload_earlySample;
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_payload = AguPlugin_setup_port_payload_earlyPc[8 : 2];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_hash = AguPlugin_setup_port_payload_pc[24 : 9];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_hit = ((Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score != 3'b000) && (Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_tag == Lsu2Plugin_logic_aguPush_0_hazardPrediction_hash));
  assign Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter = Lsu2Plugin_logic_lq_hitPrediction_mem_spinal_port1[5 : 0];
  assign Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_valid = AguPlugin_setup_port_payload_earlySample;
  assign Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_payload = AguPlugin_setup_port_payload_earlyPc[7 : 2];
  assign Lsu2Plugin_logic_aguPush_0_hitPrediction_likelyToHit = Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter[5];
  assign when_Lsu2Plugin_l733 = (Lsu2Plugin_logic_aguPush_0_pushSq && (AguPlugin_setup_port_payload_sc || AguPlugin_setup_port_payload_amo));
  assign switch_Utils_l1423_1 = AguPlugin_setup_port_payload_aguId[2:0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo = {Lsu2Plugin_logic_lq_regs_7_redo,{Lsu2Plugin_logic_lq_regs_6_redo,{Lsu2Plugin_logic_lq_regs_5_redo,{Lsu2Plugin_logic_lq_regs_4_redo,{Lsu2Plugin_logic_lq_regs_3_redo,{Lsu2Plugin_logic_lq_regs_2_redo,{Lsu2Plugin_logic_lq_regs_1_redo,Lsu2Plugin_logic_lq_regs_0_redo}}}}}}};
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo = {Lsu2Plugin_logic_sq_regs_7_redo,{Lsu2Plugin_logic_sq_regs_6_redo,{Lsu2Plugin_logic_sq_regs_5_redo,{Lsu2Plugin_logic_sq_regs_4_redo,{Lsu2Plugin_logic_sq_regs_3_redo,{Lsu2Plugin_logic_sq_regs_2_redo,{Lsu2Plugin_logic_sq_regs_1_redo,Lsu2Plugin_logic_sq_regs_0_redo}}}}}}};
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_input = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_priorityBits = Lsu2Plugin_logic_lq_ptr_priority;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask = {Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_input,(Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_input[7 : 1] & Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_priorityBits)};
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0 = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[1];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[2];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[3];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[4];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_5 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[5];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[6];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[7];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[8];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[9];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[10];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_11 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[11];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[12];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[13];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_14 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[14];
  always @(*) begin
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[0] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[1] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1 && (! Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[2] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2 && (! Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[3] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[4] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_2_to_3 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[5] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_5 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_3)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[6] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_4_to_5 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_3)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[7] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[8] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_7 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[9] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_7)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[10] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_7)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[11] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_11 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[12] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_10_to_11 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[13] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_11 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[14] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_14 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_13 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_11 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_7))));
  end

  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_2_to_3 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_3 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_4_to_5 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_5,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_4_to_5,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1}});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_7 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_7 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_7,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_4_to_5,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1}}});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_9 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_10_to_11 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_11,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_11 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_10_to_11,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_8_to_9});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_13 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pLow = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[14 : 7];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pHigh = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[6 : 0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh = (_zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh | Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pLow);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_input = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_priorityBits = Lsu2Plugin_logic_sq_ptr_priority;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask = {Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_input,(Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_input[7 : 1] & Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_priorityBits)};
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0 = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[1];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[2];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[3];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[4];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_5 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[5];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[6];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[7];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[8];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[9];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[10];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_11 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[11];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[12];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[13];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_14 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[14];
  always @(*) begin
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[0] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[1] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1 && (! Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[2] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2 && (! Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[3] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[4] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_2_to_3 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[5] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_5 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_3)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[6] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_4_to_5 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_3)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[7] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[8] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_7 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[9] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_7)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[10] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_7)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[11] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_11 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[12] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_10_to_11 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[13] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_11 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[14] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_14 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_13 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_11 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_7))));
  end

  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_2_to_3 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_3 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_4_to_5 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_5,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_4_to_5,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1}});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_7 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_7 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_7,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_4_to_5,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1}}});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_9 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_10_to_11 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_11,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_11 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_10_to_11,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_8_to_9});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_13 = (|{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12});
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pLow = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[14 : 7];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pHigh = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[6 : 0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh = (_zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh | Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pLow);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT = (|Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT = (|Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[1];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_1 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[2];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[3];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_3 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[4];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[5];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[6];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[7];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_7 = (((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_8 = (((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_1 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_9 = (((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_3 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID = {_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_9,{_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_8,_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_7}};
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[1];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_1 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[2];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[3];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_3 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[4];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[5];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[6];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[7];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_7 = (((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_8 = (((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_1 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_9 = (((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_3 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID = {_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_9,{_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_8,_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_7}};
  assign Lsu2Plugin_logic_lqSqArbitration_s0_valid = (Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT || Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ROB_FULL = {Lsu2Plugin_logic_lq_mem_robIdMsb_spinal_port1,Lsu2Plugin_logic_lq_mem_robId_spinal_port1};
  assign Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ROB_FULL = {Lsu2Plugin_logic_sq_mem_robIdMsb_spinal_port1,Lsu2Plugin_logic_sq_mem_robId_spinal_port1};
  assign Lsu2Plugin_logic_lqSqArbitration_s1_cmp = _zz_Lsu2Plugin_logic_lqSqArbitration_s1_cmp[4];
  assign Lsu2Plugin_logic_lqSqArbitration_s1_LQ_OLDER_THAN_SQ = ((! Lsu2Plugin_logic_lqSqArbitration_s1_SQ_HIT) || (Lsu2Plugin_logic_lqSqArbitration_s1_LQ_HIT && Lsu2Plugin_logic_lqSqArbitration_s1_cmp));
  assign Lsu2Plugin_logic_translationWake = Lsu2Plugin_logic_sharedPip_translationPort_wake;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION) begin
        Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_speculateHitTrapRecovered = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_sharedPip_speculateHitTrapRecovered = (Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID == 3'b000);
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION = 1'b0;
    if(when_Lsu2Plugin_l920) begin
      Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ = Lsu2Plugin_logic_lqSqArbitration_s1_LQ_OLDER_THAN_SQ;
    if(when_Lsu2Plugin_l838) begin
      Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ = 1'b0;
    end
    if(when_Lsu2Plugin_l839) begin
      Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_LQ_ROB_FULL = Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ROB_FULL;
  assign Lsu2Plugin_logic_sharedPip_stages_0_SQ_ROB_FULL = Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ROB_FULL;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_feed_takeAgu = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu[4] : _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu_1[4]);
    if(when_Lsu2Plugin_l830) begin
      Lsu2Plugin_logic_sharedPip_feed_takeAgu = 1'b1;
    end
    if(when_Lsu2Plugin_l831) begin
      Lsu2Plugin_logic_sharedPip_feed_takeAgu = 1'b0;
    end
  end

  assign when_Lsu2Plugin_l830 = (! Lsu2Plugin_logic_lqSqArbitration_s1_valid);
  assign when_Lsu2Plugin_l831 = (! AguPlugin_setup_port_valid);
  assign Lsu2Plugin_logic_sharedPip_stages_0_valid = (AguPlugin_setup_port_valid || Lsu2Plugin_logic_lqSqArbitration_s1_valid);
  assign Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l834 = (Lsu2Plugin_logic_sharedPip_feed_takeAgu || (! Lsu2Plugin_logic_sharedPip_stages_0_ready));
  assign when_Lsu2Plugin_l838 = (! Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask);
  assign when_Lsu2Plugin_l839 = (! Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask);
  assign when_Lsu2Plugin_l841 = (((Lsu2Plugin_logic_lqSqArbitration_s1_SQ_HIT && Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask) && Lsu2Plugin_logic_lqSqArbitration_s1_LQ_HIT) && Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask);
  assign Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842 = _zz_Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842;
  assign when_Lsu2Plugin_l843 = ((! Lsu2Plugin_logic_sharedPip_feed_takeAgu) && Lsu2Plugin_logic_sharedPip_stages_0_ready);
  assign when_Lsu2Plugin_l845 = (! Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ);
  assign when_Lsu2Plugin_l849 = ((Lsu2Plugin_logic_lqSqArbitration_s1_isRemoved || Lsu2Plugin_logic_lqSqArbitration_s1_ready) || (! Lsu2Plugin_logic_lqSqArbitration_s1_valid));
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID = _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID[3:0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID = _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_1[3:0];
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD = Lsu2Plugin_logic_lq_mem_physRd_spinal_port1;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD = AguPlugin_setup_port_payload_physicalRd;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_load = Lsu2Plugin_logic_lq_mem_addressPre_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_store = Lsu2Plugin_logic_sq_mem_addressPre_spinal_port1;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_load : Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_store);
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION = AguPlugin_setup_port_payload_address;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_load = Lsu2Plugin_logic_lq_mem_addressPost_spinal_port0;
  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_store = Lsu2Plugin_logic_sq_mem_addressPost_spinal_port0;
  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_load : Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_store);
  assign Lsu2Plugin_logic_sharedPip_stages_0_SIZE_load = Lsu2Plugin_logic_lq_mem_size_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_SIZE_store = Lsu2Plugin_logic_sq_mem_size_spinal_port1;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_SIZE = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_SIZE_load : Lsu2Plugin_logic_sharedPip_stages_0_SIZE_store);
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_SIZE = AguPlugin_setup_port_payload_size;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_load = Lsu2Plugin_logic_lq_mem_needTranslation_spinal_port1[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_store = Lsu2Plugin_logic_sq_mem_needTranslation_spinal_port1[0];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_load : Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_store);
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_load = Lsu2Plugin_logic_lq_mem_io_spinal_port0[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_store = Lsu2Plugin_logic_sq_mem_io_spinal_port0[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_load : Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_store);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD = Lsu2Plugin_logic_lq_mem_writeRd_spinal_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD = AguPlugin_setup_port_payload_writeRd;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_UNSIGNED = Lsu2Plugin_logic_lq_mem_unsigned_spinal_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_UNSIGNED = AguPlugin_setup_port_payload_unsigned;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LR = Lsu2Plugin_logic_lq_mem_lr_spinal_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LR = AguPlugin_setup_port_payload_lr;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC = Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port1;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC = Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port2;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID = Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_spinal_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID = Lsu2Plugin_logic_aguPush_0_hazardPrediction_hit;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA = Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_spinal_port1;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA = Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_delta;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SCORE = Lsu2Plugin_logic_lq_mem_hazardPrediction_score_spinal_port1;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SCORE = Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_AMO = Lsu2Plugin_logic_sq_mem_amo_spinal_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_AMO = AguPlugin_setup_port_payload_amo;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_SC = Lsu2Plugin_logic_sq_mem_sc_spinal_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_SC = AguPlugin_setup_port_payload_sc;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD = Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD = AguPlugin_setup_port_payload_load;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID = Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID = AguPlugin_setup_port_payload_aguId[2:0];
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID = Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID = AguPlugin_setup_port_payload_aguId[2:0];
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION_COUNTER = Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
  assign Lsu2Plugin_logic_sharedPip_stages_0_SP_FP_ADDRESS = 1'b0;
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC = AguPlugin_setup_port_payload_aguId;
  assign when_Lsu2Plugin_l920 = ((((! Lsu2Plugin_logic_lqSqArbitration_s1_valid) && AguPlugin_setup_port_payload_load) && (Lsu2Plugin_logic_aguPush_0_hitPrediction_likelyToHit || Lsu2Plugin_logic_sharedPip_stages_0_SP_FP_ADDRESS)) && Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled);
  assign Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_agu = AguPlugin_setup_port_payload_robId;
  assign Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD_agu = AguPlugin_setup_port_payload_writeRd;
  assign Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD_agu = AguPlugin_setup_port_payload_physicalRd;
  assign when_Lsu2Plugin_l929 = (AguPlugin_setup_port_valid && ((! Lsu2Plugin_logic_sharedPip_feed_takeAgu) || (! Lsu2Plugin_logic_sharedPip_stages_0_ready)));
  assign switch_Utils_l1423_2 = AguPlugin_setup_port_payload_aguId[2:0];
  assign switch_Utils_l1423_3 = AguPlugin_setup_port_payload_aguId[2:0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_isFireing = (Lsu2Plugin_logic_sharedPip_stages_0_valid && Lsu2Plugin_logic_sharedPip_stages_0_ready);
  assign Lsu2Plugin_logic_sqFeedEvent_valid = (Lsu2Plugin_logic_sharedPip_stages_0_isFireing && (! Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD));
  assign Lsu2Plugin_logic_sqFeedEvent_payload = Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID;
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = 4'bxxxx;
    case(Lsu2Plugin_logic_sharedPip_stages_0_SIZE)
      2'b00 : begin
        _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = 4'b0001;
      end
      2'b01 : begin
        _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = 4'b0011;
      end
      2'b10 : begin
        _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = (_zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK <<< Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[1 : 0]);
  assign Lsu2Plugin_logic_sharedPip_stages_0_LQCHECK_START_ID = Lsu2Plugin_logic_sq_mem_lqAlloc_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_SQCHECK_END_ID = Lsu2Plugin_logic_lq_mem_sqAlloc_spinal_port3;
  assign Lsu2Plugin_logic_sharedPip_stages_0_feed_SQ_PTR_FREE = Lsu2Plugin_logic_sq_ptr_free;
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT = (_zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT - 4'b0001);
  assign Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SQID = _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT[2:0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT = ((Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID && (! Lsu2Plugin_logic_sq_mem_feededOnce_spinal_port1[0])) && (! _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1[3]));
  assign Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_FEEDED = 1'b0;
  assign Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded = (Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED || (Lsu2Plugin_logic_sqFeedEvent_valid && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SQID)));
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded = (Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED || (Lsu2Plugin_logic_sqFeedEvent_valid && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SQID)));
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED || (Lsu2Plugin_logic_sqFeedEvent_valid && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SQID)));
  assign Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH_PC = AguPlugin_setup_port_payload_pc;
  assign when_Lsu2Plugin_l959 = (Lsu2Plugin_logic_sharedPip_stages_0_isFireing && (! Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD));
  assign Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_valid = (Lsu2Plugin_logic_sharedPip_stages_0_isFireing && Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION);
  assign Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_payload_robId = Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_agu;
  assign Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_valid = ((Lsu2Plugin_logic_sharedPip_stages_0_isFireing && Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION) && Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD_agu);
  assign Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_payload_physical = Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD_agu;
  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_valid = (|Lsu2Plugin_logic_sharedPip_stages_0_valid);
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_valid = 1'b1;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_payload_virtual = Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_payload_virtual = Lsu2Plugin_logic_special_storeAddress;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_payload_size = Lsu2Plugin_logic_sharedPip_stages_0_SIZE;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_payload_size = Lsu2Plugin_logic_special_storeSize;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_payload_redoOnDataHazard = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_payload_redoOnDataHazard = 1'b0;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_payload_unique = ((! Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD) || Lsu2Plugin_logic_sharedPip_stages_0_LR);
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_payload_unique = 1'b1;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_haltRequest_Lsu2Plugin_l990 = (! Lsu2Plugin_setup_cacheLoad_cmd_ready);
  assign when_Lsu2Plugin_l997 = (! Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION);
  always @(*) begin
    if(when_Lsu2Plugin_l997) begin
      Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_POST_TRANSLATION;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED = Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
    end
  end

  always @(*) begin
    if(when_Lsu2Plugin_l997) begin
      Lsu2Plugin_logic_sharedPip_stages_1_IS_IO = Lsu2Plugin_logic_sharedPip_stages_1_TRANSLATED_AS_IO;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_IS_IO = Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_translated_physical = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED;
    if(when_Lsu2Plugin_l1683) begin
      Lsu2Plugin_setup_cacheLoad_translated_physical = Lsu2Plugin_logic_special_storeAddress;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_translated_abord = (Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION ? ((((Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO || Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT) || Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT) || (! Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ)) || Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO) : Lsu2Plugin_logic_sharedPip_stages_1_TRANSLATED_AS_IO);
    if(when_Lsu2Plugin_l1683) begin
      Lsu2Plugin_setup_cacheLoad_translated_abord = 1'b0;
    end
  end

  assign Lsu2Plugin_setup_cacheLoad_cancels = 3'b000;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask = Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE[2 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask = {1'b0,{(3'b110 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(3'b101 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(3'b100 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(3'b011 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_1 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_2,_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_3}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID[2 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask = {1'b0,{(3'b110 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(3'b101 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(3'b100 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(3'b011 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_1 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_2,_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_3}}}}}}};
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_loopback = (Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE[3] != Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID[3]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_youngerMask = (Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_loopback ? (~ (Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask ^ Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask)) : (Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask & (~ Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask)));
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_olderMaskEmpty = (Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE == Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK = Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_youngerMask;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_NO_OLDER = Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_olderMaskEmpty;
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_pageHit = (Lsu2Plugin_logic_sq_regs_0_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_wordHit = ((Lsu2Plugin_logic_sq_regs_0_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[0] = ((((Lsu2Plugin_logic_sq_regs_0_valid && Lsu2Plugin_logic_sq_regs_0_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[0]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[1] = ((((Lsu2Plugin_logic_sq_regs_1_valid && Lsu2Plugin_logic_sq_regs_1_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[1]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[2] = ((((Lsu2Plugin_logic_sq_regs_2_valid && Lsu2Plugin_logic_sq_regs_2_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[2]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[3] = ((((Lsu2Plugin_logic_sq_regs_3_valid && Lsu2Plugin_logic_sq_regs_3_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[3]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[4] = ((((Lsu2Plugin_logic_sq_regs_4_valid && Lsu2Plugin_logic_sq_regs_4_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[4]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[5] = ((((Lsu2Plugin_logic_sq_regs_5_valid && Lsu2Plugin_logic_sq_regs_5_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[5]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[6] = ((((Lsu2Plugin_logic_sq_regs_6_valid && Lsu2Plugin_logic_sq_regs_6_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[6]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[7] = ((((Lsu2Plugin_logic_sq_regs_7_valid && Lsu2Plugin_logic_sq_regs_7_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[7]);
  end

  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_pageHit = (Lsu2Plugin_logic_sq_regs_1_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_wordHit = ((Lsu2Plugin_logic_sq_regs_1_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_pageHit = (Lsu2Plugin_logic_sq_regs_2_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_wordHit = ((Lsu2Plugin_logic_sq_regs_2_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_pageHit = (Lsu2Plugin_logic_sq_regs_3_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_wordHit = ((Lsu2Plugin_logic_sq_regs_3_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_pageHit = (Lsu2Plugin_logic_sq_regs_4_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_wordHit = ((Lsu2Plugin_logic_sq_regs_4_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_pageHit = (Lsu2Plugin_logic_sq_regs_5_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_wordHit = ((Lsu2Plugin_logic_sq_regs_5_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_pageHit = (Lsu2Plugin_logic_sq_regs_6_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_wordHit = ((Lsu2Plugin_logic_sq_regs_6_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_pageHit = (Lsu2Plugin_logic_sq_regs_7_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_wordHit = ((Lsu2Plugin_logic_sq_regs_7_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS = Lsu2Plugin_logic_sharedPip_checkSqMask_hits;
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_olderHit = ((! Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_NO_OLDER) && (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS != 8'h00));
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input = {_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[0],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[1],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[2],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[3],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[4],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[5],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[6],_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[7]}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits = Lsu2Plugin_logic_sq_ptr_priorityLast;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits = (~ {_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[0],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[1],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[2],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[3],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[4],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[5],_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[6]}}}}}});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask = {{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[6 : 0],Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[7 : 7]},(Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[6 : 0] & Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits)};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[0];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[1];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[2];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[3];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[4];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_5 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[5];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[6];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[7];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[8];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[9];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[10];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_11 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[11];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[12];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[13];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_14 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[14];
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[0] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[1] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1 && (! Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[2] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 && (! Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[3] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[4] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[5] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_5 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_3)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[6] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_3)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[7] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[8] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[9] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[10] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[11] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_11 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[12] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_10_to_11 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[13] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_11 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[14] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_14 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_11 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7))));
  end

  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_3 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_5,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1}});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1}}});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_10_to_11 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_11,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_11 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_10_to_11,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13 = (|{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pLow = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[14 : 8];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pHigh = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[7 : 0];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pHigh | _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh = {Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[0],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[1],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[2],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[3],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[4],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[5],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[6],Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[7]}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[3];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_1 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[5];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_2 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[6];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[7];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_4 = (((Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[1] || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_1) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_5 = (((Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[2] || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_2) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_6 = (((Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[4] || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_1) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_2) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel = {_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_6,{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_5,_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_4}};
  assign Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_HIT = Lsu2Plugin_logic_sharedPip_checkSqMask_olderHit;
  assign Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_ID = Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel;
  assign Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_OH = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh;
  assign Lsu2Plugin_logic_sharedPip_stages_1_isFireing = (Lsu2Plugin_logic_sharedPip_stages_1_valid && Lsu2Plugin_logic_sharedPip_stages_1_ready);
  assign when_Lsu2Plugin_l1046 = ((Lsu2Plugin_logic_sharedPip_stages_1_isFireing && Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) && (! Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT));
  assign when_Lsu2Plugin_l1052 = (Lsu2Plugin_logic_sharedPip_stages_1_isFireing && Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION);
  assign Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED = (Lsu2Plugin_logic_sq_ptr_onFreeLast_valid && (Lsu2Plugin_logic_sq_ptr_onFreeLast_payload == Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID));
  assign Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED_overloaded = ((Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED || (Lsu2Plugin_logic_sq_ptr_onFree_valid && (Lsu2Plugin_logic_sq_ptr_onFree_payload == Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID))) || ((Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID)));
  assign Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_overloaded = ((Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED || (Lsu2Plugin_logic_sq_ptr_onFree_valid && (Lsu2Plugin_logic_sq_ptr_onFree_payload == Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID))) || ((Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID)));
  assign Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_addressMatch = (Lsu2Plugin_logic_sq_mem_addressPost_spinal_port2 == Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_TRANSLATED);
  assign Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_fullMatch = ((Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_addressMatch && (Lsu2Plugin_logic_sq_mem_size_spinal_port2 == Lsu2Plugin_logic_sharedPip_stages_2_SIZE)) && (! Lsu2Plugin_logic_sq_mem_doNotBypass_spinal_port1[0]));
  assign Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_translationFailure = Lsu2Plugin_logic_sq_mem_needTranslation_spinal_port3[0];
  assign Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_data = Lsu2Plugin_logic_sq_mem_data_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_BYPASS_SUCCESS = ((! Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_translationFailure) && Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_fullMatch);
  assign Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED = Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_translationFailure;
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_endId = Lsu2Plugin_logic_lq_ptr_alloc;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask = Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID[2 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_startMask = {1'b0,{(3'b110 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(3'b101 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(3'b100 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(3'b011 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_1 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_2,_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_3}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask = Lsu2Plugin_logic_sharedPip_checkLqHits_endId[2 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_endMask = {1'b0,{(3'b110 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(3'b101 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(3'b100 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(3'b011 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_1 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_2,_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_3}}}}}}};
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_loopback = (Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID[3] != Lsu2Plugin_logic_sharedPip_checkLqHits_endId[3]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask = (Lsu2Plugin_logic_sharedPip_checkLqHits_loopback ? (~ (Lsu2Plugin_logic_sharedPip_checkLqHits_endMask ^ Lsu2Plugin_logic_sharedPip_checkLqHits_startMask)) : (Lsu2Plugin_logic_sharedPip_checkLqHits_endMask & (~ Lsu2Plugin_logic_sharedPip_checkLqHits_startMask)));
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMaskEmpty = (Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID == Lsu2Plugin_logic_sharedPip_checkLqHits_endId);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_pageHit = (Lsu2Plugin_logic_lq_regs_0_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_wordHit = ((Lsu2Plugin_logic_lq_regs_0_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_hit = ((((Lsu2Plugin_logic_lq_regs_0_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_wordHit) && Lsu2Plugin_logic_lq_regs_0_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[0]);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[0] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_hit && Lsu2Plugin_logic_lq_regs_0_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[1] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_hit && Lsu2Plugin_logic_lq_regs_1_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[2] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_hit && Lsu2Plugin_logic_lq_regs_2_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[3] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_hit && Lsu2Plugin_logic_lq_regs_3_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[4] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_hit && Lsu2Plugin_logic_lq_regs_4_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[5] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_hit && Lsu2Plugin_logic_lq_regs_5_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[6] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_hit && Lsu2Plugin_logic_lq_regs_6_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[7] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_hit && Lsu2Plugin_logic_lq_regs_7_sqChecked);
  end

  assign when_Lsu2Plugin_l1104 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_pageHit = (Lsu2Plugin_logic_lq_regs_1_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_wordHit = ((Lsu2Plugin_logic_lq_regs_1_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_hit = ((((Lsu2Plugin_logic_lq_regs_1_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_wordHit) && Lsu2Plugin_logic_lq_regs_1_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[1]);
  assign when_Lsu2Plugin_l1104_1 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_pageHit = (Lsu2Plugin_logic_lq_regs_2_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_wordHit = ((Lsu2Plugin_logic_lq_regs_2_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_hit = ((((Lsu2Plugin_logic_lq_regs_2_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_wordHit) && Lsu2Plugin_logic_lq_regs_2_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[2]);
  assign when_Lsu2Plugin_l1104_2 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_pageHit = (Lsu2Plugin_logic_lq_regs_3_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_wordHit = ((Lsu2Plugin_logic_lq_regs_3_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_hit = ((((Lsu2Plugin_logic_lq_regs_3_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_wordHit) && Lsu2Plugin_logic_lq_regs_3_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[3]);
  assign when_Lsu2Plugin_l1104_3 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_pageHit = (Lsu2Plugin_logic_lq_regs_4_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_wordHit = ((Lsu2Plugin_logic_lq_regs_4_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_hit = ((((Lsu2Plugin_logic_lq_regs_4_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_wordHit) && Lsu2Plugin_logic_lq_regs_4_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[4]);
  assign when_Lsu2Plugin_l1104_4 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_pageHit = (Lsu2Plugin_logic_lq_regs_5_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_wordHit = ((Lsu2Plugin_logic_lq_regs_5_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_hit = ((((Lsu2Plugin_logic_lq_regs_5_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_wordHit) && Lsu2Plugin_logic_lq_regs_5_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[5]);
  assign when_Lsu2Plugin_l1104_5 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_pageHit = (Lsu2Plugin_logic_lq_regs_6_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_wordHit = ((Lsu2Plugin_logic_lq_regs_6_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_hit = ((((Lsu2Plugin_logic_lq_regs_6_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_wordHit) && Lsu2Plugin_logic_lq_regs_6_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[6]);
  assign when_Lsu2Plugin_l1104_6 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_pageHit = (Lsu2Plugin_logic_lq_regs_7_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_wordHit = ((Lsu2Plugin_logic_lq_regs_7_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_hit = ((((Lsu2Plugin_logic_lq_regs_7_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_wordHit) && Lsu2Plugin_logic_lq_regs_7_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[7]);
  assign when_Lsu2Plugin_l1104_7 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_hit);
  assign Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER = Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMaskEmpty;
  assign Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerHit = ((Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS != 8'h00) && (! Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_NO_YOUNGER));
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_input = Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_priorityBits = Lsu2Plugin_logic_lq_ptr_priorityLast;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask = {Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_input,(Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_input[7 : 1] & Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_priorityBits)};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 = Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[0];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[1];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[2];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[3];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[4];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_5 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[5];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[6];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[7];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[8];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[9];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[10];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_11 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[11];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[12];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[13];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_14 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[14];
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[0] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[1] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1 && (! Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[2] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 && (! Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[3] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[4] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[5] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_5 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_3)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[6] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_3)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[7] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[8] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[9] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[10] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[11] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_11 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[12] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_10_to_11 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[13] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_11 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[14] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_14 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_11 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7))));
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_3 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_5,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1}});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_7 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_4_to_5,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_2_to_3,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1}}});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_10_to_11 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_11,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_11 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_10_to_11,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_8_to_9});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13 = (|{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12});
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pLow = Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[14 : 7];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pHigh = Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[6 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh = (_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh | Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pLow);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[3];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_1 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[5];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_2 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[6];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[7];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_4 = (((Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[1] || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_1) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_5 = (((Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[2] || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_2) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_6 = (((Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[4] || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_1) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_2) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3);
  assign Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel = {_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_6,{_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_5,_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_4}};
  assign Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ROB = Lsu2Plugin_logic_lq_mem_robId_spinal_port2;
  assign Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_RESCHEDULE = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerHit;
  assign Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ID = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride = 1'b1;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride = 1'b1;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_valid = Lsu2Plugin_setup_cacheLoad_rsp_valid;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data = Lsu2Plugin_setup_cacheLoad_rsp_payload_data;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data = LsuPlugin_peripheralBus_rsp_payload_data;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_fault = Lsu2Plugin_setup_cacheLoad_rsp_payload_fault;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_redo = Lsu2Plugin_setup_cacheLoad_rsp_payload_redo;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlot = Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlot;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlotAny = Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlotAny;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize = Lsu2Plugin_logic_sharedPip_stages_2_SIZE;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize = Lsu2Plugin_logic_special_loadSize;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize = Lsu2Plugin_logic_special_storeSize;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress = Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress = Lsu2Plugin_logic_special_loadAddress;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress = Lsu2Plugin_logic_special_storeAddress;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned = Lsu2Plugin_logic_sharedPip_stages_2_UNSIGNED;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned = Lsu2Plugin_logic_special_loadUnsigned;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_0 = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data[7 : 0];
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_1 = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data[15 : 8];
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_2 = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data[23 : 16];
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3 = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data[31 : 24];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[7 : 0] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted;
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[15 : 8] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_2;
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[23 : 16] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_2;
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[31 : 24] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3;
    if(when_Lsu2Plugin_l1158) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_data;
    end
  end

  assign when_Lsu2Plugin_l1158 = ((! Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride) && Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_HIT);
  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = (Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[7] && (! Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned));
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[31] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[30] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[29] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[28] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[27] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[26] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[25] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[24] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[23] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[22] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[21] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[20] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[19] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[18] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[17] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[16] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[15] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[14] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[13] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[12] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[11] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[10] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[9] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[8] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[7 : 0] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[7 : 0];
  end

  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2 = (Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[15] && (! Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned));
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[31] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[30] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[29] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[28] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[27] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[26] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[25] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[24] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[23] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[22] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[21] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[20] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[19] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[18] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[17] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[16] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[15 : 0] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[15 : 0];
  end

  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_4[31 : 0] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[31 : 0];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize)
      2'b00 : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1;
      end
      2'b01 : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3;
      end
      2'b10 : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_4;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_isFireing = (Lsu2Plugin_logic_sharedPip_stages_2_valid && Lsu2Plugin_logic_sharedPip_stages_2_ready);
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_valid = ((Lsu2Plugin_logic_sharedPip_stages_2_isFireing && (! Lsu2Plugin_logic_sharedPip_stages_2_IS_IO)) && ((! Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION) || ((! Lsu2Plugin_logic_sharedPip_stages_2_MMU_REDO) && (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT))));
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_isLoad = Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_address = Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_TRANSLATED;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_readData = Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_robId = Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_lqId = Lsu2Plugin_logic_sharedPip_stages_2_LQ_ID;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_size = Lsu2Plugin_logic_sharedPip_stages_2_SIZE;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_doIt = (((Lsu2Plugin_logic_sharedPip_stages_2_valid && Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD) && Lsu2Plugin_logic_sharedPip_stages_2_WRITE_RD) && ((! Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION) || ((Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_READ && (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT)) && (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_ACCESS_FAULT))));
  always @(*) begin
    Lsu2Plugin_setup_regfilePorts_0_write_valid = ((Lsu2Plugin_logic_sharedPip_cacheRsp_doIt && Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD) && 1'b1);
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_regfilePorts_0_write_valid = (Lsu2Plugin_logic_special_loadWriteRd && 1'b1);
    end
    if(Lsu2Plugin_logic_special_atomic_comp_rfWrite) begin
      Lsu2Plugin_setup_regfilePorts_0_write_valid = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_regfilePorts_0_write_address = Lsu2Plugin_logic_sharedPip_stages_2_PHYS_RD;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_regfilePorts_0_write_address = Lsu2Plugin_logic_special_loadPhysRd;
    end
    if(Lsu2Plugin_logic_special_atomic_comp_rfWrite) begin
      Lsu2Plugin_setup_regfilePorts_0_write_address = Lsu2Plugin_logic_sq_mem_physRd;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_regfilePorts_0_write_data = Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
        Lsu2Plugin_setup_regfilePorts_0_write_data = 32'h00000000;
        Lsu2Plugin_setup_regfilePorts_0_write_data[0] = (! Lsu2Plugin_logic_special_atomic_gotReservation);
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_regfilePorts_0_write_robId = Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_regfilePorts_0_write_robId = Lsu2Plugin_logic_special_robId;
    end
    if(Lsu2Plugin_logic_special_atomic_comp_rfWrite) begin
      Lsu2Plugin_setup_regfilePorts_0_write_robId = Lsu2Plugin_logic_special_robId;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_fpuWriteSize = Lsu2Plugin_logic_sharedPip_stages_2_SIZE;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_fpuWriteSize = Lsu2Plugin_logic_special_loadSize;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_WRITE_FAILURE = ((Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride) && (! Lsu2Plugin_logic_sharedPip_stages_2_IS_IO));
  assign Lsu2Plugin_logic_sharedPip_stages_2_MISS_ALIGNED = (|{((Lsu2Plugin_logic_sharedPip_stages_2_SIZE == 2'b10) && (Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION[1 : 0] != 2'b00)),((Lsu2Plugin_logic_sharedPip_stages_2_SIZE == 2'b01) && (Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION[0 : 0] != 1'b0))});
  assign Lsu2Plugin_logic_sharedPip_stages_2_PAGE_FAULT = ((Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD ? (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_READ) : (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_WRITE)) || Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_success = 1'b0;
    if(!Lsu2Plugin_logic_sharedPip_stages_2_MISS_ALIGNED) begin
      if(!when_Lsu2Plugin_l1203) begin
        if(!when_Lsu2Plugin_l1205) begin
          if(!when_Lsu2Plugin_l1207) begin
            if(!when_Lsu2Plugin_l1209) begin
              if(!when_Lsu2Plugin_l1211) begin
                if(!when_Lsu2Plugin_l1213) begin
                  Lsu2Plugin_logic_sharedPip_cacheRsp_success = 1'b1;
                end
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_stages_2_MISS_ALIGNED) begin
      Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN;
    end else begin
      if(when_Lsu2Plugin_l1203) begin
        Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_MMU_REDO;
      end else begin
        if(when_Lsu2Plugin_l1205) begin
          Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_TRAP_MMU;
        end else begin
          if(when_Lsu2Plugin_l1207) begin
            Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD;
          end else begin
            if(when_Lsu2Plugin_l1209) begin
              Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_LOAD_MISS;
            end else begin
              if(when_Lsu2Plugin_l1211) begin
                Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_LOAD_FAILED;
              end else begin
                if(when_Lsu2Plugin_l1213) begin
                  Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS;
                end else begin
                  Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_SUCCESS;
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_Lsu2Plugin_l1203 = (Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION && Lsu2Plugin_logic_sharedPip_stages_2_MMU_REDO);
  assign when_Lsu2Plugin_l1205 = (Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION && (Lsu2Plugin_logic_sharedPip_stages_2_MMU_ACCESS_FAULT || Lsu2Plugin_logic_sharedPip_stages_2_PAGE_FAULT));
  assign when_Lsu2Plugin_l1207 = (Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && ((Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_HIT && (! Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_BYPASS_SUCCESS)) || Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT));
  assign when_Lsu2Plugin_l1209 = (Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_redo);
  assign when_Lsu2Plugin_l1211 = (Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && Lsu2Plugin_logic_sharedPip_stages_2_LOAD_WRITE_FAILURE);
  assign when_Lsu2Plugin_l1213 = (Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_fault);
  assign Lsu2Plugin_logic_sharedPip_stages_2_TRAP_SPECULATION = (Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION && ((! Lsu2Plugin_logic_sharedPip_cacheRsp_success) || Lsu2Plugin_logic_sharedPip_stages_2_IS_IO));
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_valid = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_data = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_fault = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_fault;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_redo = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_redo;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny = (Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlotAny && (! (|DataCachePlugin_setup_refillCompletions)));
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlot = (Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlot & (~ DataCachePlugin_setup_refillCompletions));
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_valid = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_data = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_data;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_fault = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_fault;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_redo = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_redo;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlotAny && (! (|DataCachePlugin_setup_refillCompletions)));
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlot = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlot & (~ DataCachePlugin_setup_refillCompletions));
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC = (Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD ? Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID : Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ID);
  assign Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC = Lsu2Plugin_logic_lq_mem_pc_spinal_port1;
  always @(*) begin
    Lsu2Plugin_setup_sharedCompletion_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(when_Lsu2Plugin_l1333) begin
              Lsu2Plugin_setup_sharedCompletion_valid = 1'b1;
            end
          end else begin
            if(when_Lsu2Plugin_l1374) begin
              Lsu2Plugin_setup_sharedCompletion_valid = 1'b1;
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_setup_sharedCompletion_payload_id = Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(when_Lsu2Plugin_l1333) begin
              if(when_Lsu2Plugin_l1335) begin
                Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_valid = 1'b1;
              end
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_payload_robId = Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(when_Lsu2Plugin_l1333) begin
              if(when_Lsu2Plugin_l1335) begin
                Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid = 1'b1;
              end
            end
          end
        end
      endcase
    end
    if(Lsu2Plugin_logic_special_atomic_comp_wakeRf) begin
      Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_payload_physical = Lsu2Plugin_logic_sharedPip_stages_3_PHYS_RD;
    if(Lsu2Plugin_logic_special_atomic_comp_wakeRf) begin
      Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_payload_physical = Lsu2Plugin_logic_sq_mem_physRd;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION) begin
        Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
      end
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
          Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
          Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
          Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_payload_robId = Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_setup_sharedTrap_payload_robId = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ROB;
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_setup_sharedTrap_payload_tval = Lsu2Plugin_logic_sharedPip_stages_3_ADDRESS_PRE_TRANSLATION;
  assign Lsu2Plugin_setup_sharedTrap_payload_skipCommit = 1'b1;
  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_payload_trap = 1'b1;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_setup_sharedTrap_payload_trap = 1'b0;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_payload_cause = 4'bxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION) begin
        Lsu2Plugin_setup_sharedTrap_payload_cause = 4'b1010;
      end
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
          Lsu2Plugin_setup_sharedTrap_payload_cause = 4'b0100;
          Lsu2Plugin_setup_sharedTrap_payload_cause[1] = (! Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD);
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
          Lsu2Plugin_setup_sharedTrap_payload_cause = 4'b1101;
          Lsu2Plugin_setup_sharedTrap_payload_cause[1] = (! Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD);
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
          Lsu2Plugin_setup_sharedTrap_payload_cause = 4'b0101;
          Lsu2Plugin_setup_sharedTrap_payload_cause[1] = (! Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_payload_reason = 8'bxxxxxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION) begin
        Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h03;
      end
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
          Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h01;
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
          Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h01;
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
          Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h01;
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h20;
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_setup_sharedTrap_payload_pcTarget = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC;
  assign Lsu2Plugin_logic_sharedPip_ctrl_lqMask = (8'h01 <<< Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID);
  assign Lsu2Plugin_logic_sharedPip_ctrl_sqMask = (8'h01 <<< Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger = Lsu2Plugin_logic_translationWake;
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger = (! (|Lsu2Plugin_logic_sharedPip_ctrl_refillMask));
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
          Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger = 1'b1;
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign _zz_118 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[0];
  assign _zz_119 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[1];
  assign _zz_120 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[2];
  assign _zz_121 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[3];
  assign _zz_122 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[4];
  assign _zz_123 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[5];
  assign _zz_124 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[6];
  assign _zz_125 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[7];
  assign _zz_126 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[0];
  assign _zz_127 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[1];
  assign _zz_128 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[2];
  assign _zz_129 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[3];
  assign _zz_130 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[4];
  assign _zz_131 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[5];
  assign _zz_132 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[6];
  assign _zz_133 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[7];
  assign Lsu2Plugin_logic_sharedPip_ctrl_refillMask = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlotAny ? 2'b11 : Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlot);
  assign Lsu2Plugin_logic_sharedPip_ctrl_doCompletion = ((Lsu2Plugin_logic_sharedPip_stages_3_CTRL == Lsu2Plugin_CTRL_ENUM_SUCCESS) && (! Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION));
  assign Lsu2Plugin_logic_sharedPip_stages_3_isFireing = (Lsu2Plugin_logic_sharedPip_stages_3_valid && Lsu2Plugin_logic_sharedPip_stages_3_ready);
  assign when_Lsu2Plugin_l1313 = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT || Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_WAIT_FEED);
  assign _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT ? Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SQID : Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID);
  assign when_Lsu2Plugin_l1314 = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT ? Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_resulting : Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_resulting);
  assign when_Lsu2Plugin_l1333 = (! Lsu2Plugin_logic_sharedPip_stages_3_IS_IO);
  assign when_Lsu2Plugin_l1335 = (Lsu2Plugin_logic_sharedPip_stages_3_WRITE_RD && (! Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION));
  assign _zz_when_Lsu2Plugin_l1348 = _zz__zz_when_Lsu2Plugin_l1348;
  always @(*) begin
    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'b000;
    if(when_Lsu2Plugin_l1348) begin
      _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'b001;
    end
    if(when_Lsu2Plugin_l1351) begin
      _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'b111;
    end
  end

  assign when_Lsu2Plugin_l1348 = (_zz_when_Lsu2Plugin_l1348 && (&Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE));
  assign when_Lsu2Plugin_l1351 = ((! _zz_when_Lsu2Plugin_l1348) && (! (|Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE)));
  assign when_Lsu2Plugin_l1374 = (((! Lsu2Plugin_logic_sharedPip_stages_3_SC) && (! Lsu2Plugin_logic_sharedPip_stages_3_AMO)) && (! Lsu2Plugin_logic_sharedPip_stages_3_IS_IO));
  assign _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next = ((Lsu2Plugin_logic_sharedPip_ctrl_doCompletion && (! Lsu2Plugin_logic_sharedPip_stages_3_IS_IO)) ? 6'h3f : 6'h14);
  assign Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next = ($signed(_zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_1) + $signed(_zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_2));
  assign Lsu2Plugin_logic_lq_hitPrediction_write_valid = (((Lsu2Plugin_logic_sharedPip_stages_3_isFireing && Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) && Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH) && (! Lsu2Plugin_logic_sharedPip_stages_3_SP_FP_ADDRESS));
  assign Lsu2Plugin_logic_lq_hitPrediction_write_payload_address = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH_PC[7 : 2];
  assign when_SInt_l131 = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[6];
  assign when_SInt_l132 = (! (&_zz_when_SInt_l132));
  always @(*) begin
    if(when_SInt_l131) begin
      if(when_SInt_l132) begin
        _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = 6'h20;
      end else begin
        _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[5 : 0];
      end
    end else begin
      if(when_SInt_l138) begin
        _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = 6'h1f;
      end else begin
        _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[5 : 0];
      end
    end
  end

  assign when_SInt_l138 = (|_zz_when_SInt_l138);
  assign Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter;
  assign Lsu2Plugin_logic_writeback_waitOn_ready = ((Lsu2Plugin_logic_writeback_waitOn_refillSlot == 2'b00) && (! Lsu2Plugin_logic_writeback_waitOn_refillSlotAny));
  always @(*) begin
    Lsu2Plugin_logic_writeback_waitOn_refillSlotSet = 2'b00;
    if(when_Lsu2Plugin_l1488) begin
      if(Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        Lsu2Plugin_logic_writeback_waitOn_refillSlotSet = Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlot;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_writeback_waitOn_refillSlotAnySet = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      if(Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        Lsu2Plugin_logic_writeback_waitOn_refillSlotAnySet = Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlotAny;
      end
    end
  end

  assign Lsu2Plugin_logic_writeback_feed_holdPrefetch = 1'b0;
  always @(*) begin
    Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready = toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready;
    if(when_Stream_l369_2) begin
      Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l369_2 = (! toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_valid);
  assign toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_valid = toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rValid;
  assign toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_payload = toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rData;
  assign _zz_toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready = (! Lsu2Plugin_logic_writeback_feed_holdPrefetch);
  assign toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready = (1'b1 && _zz_toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready);
  assign Lsu2Plugin_logic_writeback_feed_prediction_valid = (toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_valid && _zz_toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready);
  assign Lsu2Plugin_logic_writeback_feed_prediction_payload = toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_payload;
  assign Lsu2Plugin_logic_writeback_feed_io = Lsu2Plugin_logic_sq_mem_io_spinal_port2[0];
  assign Lsu2Plugin_logic_writeback_feed_size = Lsu2Plugin_logic_sq_mem_size_spinal_port3;
  always @(*) begin
    Lsu2Plugin_logic_writeback_feed_data = Lsu2Plugin_logic_sq_mem_data_spinal_port2;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
        if(Lsu2Plugin_logic_special_storeAmo) begin
          Lsu2Plugin_logic_writeback_feed_data[31 : 0] = Lsu2Plugin_logic_special_atomic_result;
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_logic_writeback_feed_skip = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
        if(when_Lsu2Plugin_l1828) begin
          Lsu2Plugin_logic_writeback_feed_skip = 1'b1;
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_writeback_feed_doit = (((Lsu2Plugin_logic_sq_ptr_writeBack != Lsu2Plugin_logic_sq_ptr_commit) && Lsu2Plugin_logic_writeback_waitOn_ready) && (! Lsu2Plugin_logic_writeback_feed_prediction_valid));
  always @(*) begin
    Lsu2Plugin_logic_writeback_feed_fire = (Lsu2Plugin_logic_writeback_feed_doit && Lsu2Plugin_setup_cacheStore_cmd_ready);
    if(when_Lsu2Plugin_l1509) begin
      Lsu2Plugin_logic_writeback_feed_fire = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_valid = Lsu2Plugin_logic_writeback_feed_doit;
    if(Lsu2Plugin_logic_writeback_feed_prediction_valid) begin
      Lsu2Plugin_setup_cacheStore_cmd_valid = 1'b1;
    end
    if(when_Lsu2Plugin_l1509) begin
      Lsu2Plugin_setup_cacheStore_cmd_valid = 1'b0;
    end
    if(when_Lsu2Plugin_l1553) begin
      Lsu2Plugin_setup_cacheStore_cmd_valid = (! Lsu2Plugin_logic_flush_cmdPtr[2]);
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_address = Lsu2Plugin_logic_sq_mem_addressPost_spinal_port3;
    if(Lsu2Plugin_logic_writeback_feed_prediction_valid) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_address = Lsu2Plugin_logic_writeback_feed_prediction_payload;
    end
    if(when_Lsu2Plugin_l1553) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_address[7 : 6] = Lsu2Plugin_logic_flush_cmdPtr[1:0];
    end
  end

  always @(*) begin
    _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask = 4'bxxxx;
    case(Lsu2Plugin_logic_writeback_feed_size)
      2'b00 : begin
        _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask = 4'b0001;
      end
      2'b01 : begin
        _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask = 4'b0011;
      end
      2'b10 : begin
        _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_cacheStore_cmd_payload_mask = (_zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask <<< Lsu2Plugin_setup_cacheStore_cmd_payload_address[1 : 0]);
  assign Lsu2Plugin_setup_cacheStore_cmd_payload_generation = Lsu2Plugin_logic_writeback_generation;
  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(Lsu2Plugin_logic_writeback_feed_size)
      2'b00 : begin
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[7 : 0] = Lsu2Plugin_logic_writeback_feed_data[7 : 0];
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[15 : 8] = Lsu2Plugin_logic_writeback_feed_data[7 : 0];
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[23 : 16] = Lsu2Plugin_logic_writeback_feed_data[7 : 0];
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[31 : 24] = Lsu2Plugin_logic_writeback_feed_data[7 : 0];
      end
      2'b01 : begin
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[15 : 0] = Lsu2Plugin_logic_writeback_feed_data[15 : 0];
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[31 : 16] = Lsu2Plugin_logic_writeback_feed_data[15 : 0];
      end
      2'b10 : begin
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[31 : 0] = Lsu2Plugin_logic_writeback_feed_data[31 : 0];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_io = Lsu2Plugin_logic_writeback_feed_io;
    if(Lsu2Plugin_logic_writeback_feed_prediction_valid) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_io = 1'b0;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_prefetch = 1'b0;
    if(Lsu2Plugin_logic_writeback_feed_prediction_valid) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_prefetch = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_valid = Lsu2Plugin_setup_cacheStore_rsp_valid;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_fault = Lsu2Plugin_setup_cacheStore_rsp_payload_fault;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_redo = Lsu2Plugin_setup_cacheStore_rsp_payload_redo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlot = Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlot;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlotAny = Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlotAny;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_generationKo = Lsu2Plugin_setup_cacheStore_rsp_payload_generationKo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_flush = Lsu2Plugin_setup_cacheStore_rsp_payload_flush;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_prefetch = Lsu2Plugin_setup_cacheStore_rsp_payload_prefetch;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_address = Lsu2Plugin_setup_cacheStore_rsp_payload_address;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_io = Lsu2Plugin_setup_cacheStore_rsp_payload_io;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_valid = Lsu2Plugin_logic_writeback_rsp_delayed_0_valid;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_fault = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_fault;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_redo = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_redo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_generationKo = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_generationKo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_flush = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_flush;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_prefetch = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_prefetch;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_address = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_address;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_io = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_io;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_valid = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_valid;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_fault = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_fault;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_redo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlot = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlot;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlotAny = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlotAny;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_generationKo = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_generationKo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_flush = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_flush;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_prefetch = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_prefetch;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_address = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_address;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_io = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_io;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlot = (Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlot & (~ DataCachePlugin_setup_refillCompletions));
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlotAny = (Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlotAny && (DataCachePlugin_setup_refillCompletions == 2'b00));
  always @(*) begin
    Lsu2Plugin_logic_sq_ptr_onFree_valid = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      if(!Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        Lsu2Plugin_logic_sq_ptr_onFree_valid = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l1509) begin
      Lsu2Plugin_logic_sq_ptr_onFree_valid = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_sq_ptr_onFree_payload = Lsu2Plugin_logic_sq_ptr_freeReal;
  always @(*) begin
    Lsu2Plugin_logic_writeback_rsp_whitebox_valid = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      if(!Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        if(when_Lsu2Plugin_l1498) begin
          Lsu2Plugin_logic_writeback_rsp_whitebox_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_prefetch_predictor_io_learn_valid = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      Lsu2Plugin_logic_prefetch_predictor_io_learn_valid = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_prefetch_predictor_io_learn_payload_allocate = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      if(Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        Lsu2Plugin_logic_prefetch_predictor_io_learn_payload_allocate = 1'b1;
      end
    end
  end

  assign when_Lsu2Plugin_l1488 = (((Lsu2Plugin_logic_writeback_rsp_delayed_1_valid && (! Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_generationKo)) && (! Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_flush)) && (! Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_prefetch));
  assign when_Lsu2Plugin_l1498 = (! Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_io);
  assign Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_valid = (Lsu2Plugin_logic_writeback_rsp_delayed_1_valid && Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_prefetch);
  assign Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_payload = (|Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlot);
  assign when_Lsu2Plugin_l1509 = (Lsu2Plugin_logic_writeback_feed_doit && Lsu2Plugin_logic_writeback_feed_skip);
  always @(*) begin
    Lsu2Plugin_logic_sq_tracker_add = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      Lsu2Plugin_logic_sq_tracker_add = 1'b1;
    end
  end

  assign when_Lsu2Plugin_l1521 = (Lsu2Plugin_logic_sq_ptr_priority == 7'h00);
  assign when_Lsu2Plugin_l1524 = (Lsu2Plugin_logic_sq_ptr_freeReal == 3'b000);
  assign when_Lsu2Plugin_l1524_1 = (Lsu2Plugin_logic_sq_ptr_freeReal == 3'b001);
  assign when_Lsu2Plugin_l1524_2 = (Lsu2Plugin_logic_sq_ptr_freeReal == 3'b010);
  assign when_Lsu2Plugin_l1524_3 = (Lsu2Plugin_logic_sq_ptr_freeReal == 3'b011);
  assign when_Lsu2Plugin_l1524_4 = (Lsu2Plugin_logic_sq_ptr_freeReal == 3'b100);
  assign when_Lsu2Plugin_l1524_5 = (Lsu2Plugin_logic_sq_ptr_freeReal == 3'b101);
  assign when_Lsu2Plugin_l1524_6 = (Lsu2Plugin_logic_sq_ptr_freeReal == 3'b110);
  assign when_Lsu2Plugin_l1524_7 = (Lsu2Plugin_logic_sq_ptr_freeReal == 3'b111);
  assign FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548 = _zz_FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548;
  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_flush = 1'b0;
    if(when_Lsu2Plugin_l1553) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_flush = 1'b1;
    end
  end

  assign Lsu2Plugin_setup_cacheStore_cmd_payload_flushFree = Lsu2Plugin_logic_flush_withFree;
  assign when_Lsu2Plugin_l1553 = (Lsu2Plugin_logic_flush_busy && Lsu2Plugin_logic_flush_doit);
  assign Lsu2Plugin_setup_cacheStore_cmd_fire = (Lsu2Plugin_setup_cacheStore_cmd_valid && Lsu2Plugin_setup_cacheStore_cmd_ready);
  assign when_Lsu2Plugin_l1561 = (Lsu2Plugin_setup_cacheStore_rsp_valid && (! Lsu2Plugin_setup_cacheStore_rsp_payload_generationKo));
  assign when_Lsu2Plugin_l1569 = (Lsu2Plugin_logic_flush_rspPtr[2] && (! DataCachePlugin_setup_writebackBusy));
  assign Lsu2Plugin_logic_special_lqOnTop = (Lsu2Plugin_logic_lq_mem_robId_spinal_port3 == CommitPlugin_logic_commit_head);
  assign Lsu2Plugin_logic_special_sqOnTop = (Lsu2Plugin_logic_sq_mem_robId_spinal_port2 == CommitPlugin_logic_commit_head);
  assign Lsu2Plugin_logic_special_storeWriteBackUsable = (Lsu2Plugin_logic_sq_ptr_writeBack == Lsu2Plugin_logic_sq_ptr_commit);
  assign Lsu2Plugin_logic_special_storeSpecial = Lsu2Plugin_logic_sq_mem_doSpecial_spinal_port2[0];
  assign Lsu2Plugin_logic_special_loadSpecial = Lsu2Plugin_logic_lq_mem_doSpecial_spinal_port2[0];
  assign Lsu2Plugin_logic_special_storeHit = (((Lsu2Plugin_logic_special_sqOnTop && Lsu2Plugin_logic_special_storeWriteBackUsable) && (Lsu2Plugin_logic_sq_ptr_commit != Lsu2Plugin_logic_sq_ptr_alloc)) && Lsu2Plugin_logic_special_storeSpecial);
  assign Lsu2Plugin_logic_special_loadHit = ((Lsu2Plugin_logic_special_lqOnTop && (Lsu2Plugin_logic_lq_ptr_free != Lsu2Plugin_logic_lq_ptr_alloc)) && Lsu2Plugin_logic_special_loadSpecial);
  assign Lsu2Plugin_logic_special_hit = (Lsu2Plugin_logic_special_storeHit || Lsu2Plugin_logic_special_loadHit);
  always @(*) begin
    Lsu2Plugin_logic_special_fire = LsuPlugin_peripheralBus_rsp_valid_regNext;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
        if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
          Lsu2Plugin_logic_special_fire = 1'b1;
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign LsuPlugin_peripheralBus_cmd_fire = (LsuPlugin_peripheralBus_cmd_valid && LsuPlugin_peripheralBus_cmd_ready);
  assign Lsu2Plugin_logic_special_address = (Lsu2Plugin_logic_special_isStore ? Lsu2Plugin_logic_special_storeAddress : Lsu2Plugin_logic_special_loadAddress);
  assign Lsu2Plugin_logic_special_addressVirt = (Lsu2Plugin_logic_special_isStore ? Lsu2Plugin_logic_special_storeAddressVirt : Lsu2Plugin_logic_special_loadAddressVirt);
  assign Lsu2Plugin_logic_special_isIo = (! (Lsu2Plugin_logic_special_isStore && (Lsu2Plugin_logic_special_storeAmo || Lsu2Plugin_logic_special_storeSc)));
  assign Lsu2Plugin_logic_special_isAtomic = (! Lsu2Plugin_logic_special_isIo);
  always @(*) begin
    Lsu2Plugin_logic_special_wakeRob_valid = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      if(Lsu2Plugin_logic_special_loadWriteRd) begin
        Lsu2Plugin_logic_special_wakeRob_valid = 1'b1;
      end
    end
    if(Lsu2Plugin_logic_special_atomic_comp_wakeRf) begin
      Lsu2Plugin_logic_special_wakeRob_valid = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_special_wakeRob_payload_robId = Lsu2Plugin_logic_special_robId;
  always @(*) begin
    Lsu2Plugin_logic_special_wakeRf_valid = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      if(Lsu2Plugin_logic_special_loadWriteRd) begin
        Lsu2Plugin_logic_special_wakeRf_valid = 1'b1;
      end
    end
  end

  assign Lsu2Plugin_logic_special_wakeRf_payload_physical = Lsu2Plugin_logic_special_loadPhysRd;
  assign LsuPlugin_peripheralBus_cmd_valid = ((Lsu2Plugin_logic_special_enabled && (! Lsu2Plugin_logic_special_cmdSent)) && Lsu2Plugin_logic_special_isIo);
  assign LsuPlugin_peripheralBus_cmd_payload_write = Lsu2Plugin_logic_special_isStore;
  assign LsuPlugin_peripheralBus_cmd_payload_address = Lsu2Plugin_logic_special_address;
  assign LsuPlugin_peripheralBus_cmd_payload_size = (Lsu2Plugin_logic_special_isStore ? Lsu2Plugin_logic_special_storeSize : Lsu2Plugin_logic_special_loadSize);
  assign LsuPlugin_peripheralBus_cmd_payload_data = Lsu2Plugin_logic_special_storeData;
  assign LsuPlugin_peripheralBus_cmd_payload_mask = Lsu2Plugin_logic_special_storeMask;
  always @(*) begin
    Lsu2Plugin_setup_specialTrap_valid = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_specialTrap_valid = LsuPlugin_peripheralBus_rsp_payload_error;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
        Lsu2Plugin_setup_specialTrap_valid = 1'b1;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_specialTrap_payload_robId = Lsu2Plugin_logic_special_robId;
  assign Lsu2Plugin_setup_specialTrap_payload_cause = {1'd0, _zz_Lsu2Plugin_setup_specialTrap_payload_cause};
  assign Lsu2Plugin_setup_specialTrap_payload_tval = Lsu2Plugin_logic_special_addressVirt;
  assign Lsu2Plugin_setup_specialTrap_payload_skipCommit = 1'b1;
  assign Lsu2Plugin_setup_specialTrap_payload_reason = 8'h01;
  always @(*) begin
    Lsu2Plugin_setup_specialCompletion_valid = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_specialCompletion_valid = 1'b1;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
        Lsu2Plugin_setup_specialCompletion_valid = 1'b1;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_specialCompletion_payload_id = Lsu2Plugin_logic_special_robId;
  assign Lsu2Plugin_logic_special_atomic_wantExit = 1'b0;
  always @(*) begin
    Lsu2Plugin_logic_special_atomic_wantStart = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
        Lsu2Plugin_logic_special_atomic_wantStart = 1'b1;
      end
    endcase
  end

  assign Lsu2Plugin_logic_special_atomic_wantKill = 1'b0;
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub = Lsu2Plugin_logic_special_atomic_readed[31 : 0];
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 = Lsu2Plugin_logic_special_storeData[31 : 0];
  assign Lsu2Plugin_logic_special_atomic_alu_compare = Lsu2Plugin_logic_sq_mem_op[2];
  assign Lsu2Plugin_logic_special_atomic_alu_unsigned = Lsu2Plugin_logic_sq_mem_op[1];
  assign Lsu2Plugin_logic_special_atomic_alu_addSub = _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_2;
  assign Lsu2Plugin_logic_special_atomic_alu_less = ((_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1[31] == _zz_Lsu2Plugin_logic_special_atomic_alu_addSub[31]) ? Lsu2Plugin_logic_special_atomic_alu_addSub[31] : (Lsu2Plugin_logic_special_atomic_alu_unsigned ? _zz_Lsu2Plugin_logic_special_atomic_alu_addSub[31] : _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1[31]));
  assign Lsu2Plugin_logic_special_atomic_alu_selectRf = (Lsu2Plugin_logic_sq_mem_swap ? 1'b1 : (Lsu2Plugin_logic_sq_mem_op[0] ^ Lsu2Plugin_logic_special_atomic_alu_less));
  assign switch_Misc_l241_1 = (Lsu2Plugin_logic_sq_mem_op | {Lsu2Plugin_logic_sq_mem_swap,2'b00});
  always @(*) begin
    case(switch_Misc_l241_1)
      3'b000 : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = Lsu2Plugin_logic_special_atomic_alu_addSub;
      end
      3'b001 : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = (_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 ^ _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
      end
      3'b010 : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = (_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 | _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
      end
      3'b011 : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = (_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 & _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
      end
      default : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = (Lsu2Plugin_logic_special_atomic_alu_selectRf ? _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 : _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
      end
    endcase
  end

  assign Lsu2Plugin_logic_special_atomic_alu_result = Lsu2Plugin_logic_special_atomic_alu_raw;
  assign when_Lsu2Plugin_l1683 = (Lsu2Plugin_logic_special_enabled && Lsu2Plugin_logic_special_isAtomic);
  always @(*) begin
    DataCachePlugin_setup_lockPort_valid = 1'b0;
    if(when_Lsu2Plugin_l1698) begin
      DataCachePlugin_setup_lockPort_valid = 1'b1;
    end
  end

  always @(*) begin
    DataCachePlugin_setup_lockPort_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_Lsu2Plugin_l1698) begin
      DataCachePlugin_setup_lockPort_address = Lsu2Plugin_logic_special_storeAddress;
    end
  end

  assign Lsu2Plugin_setup_cacheLoad_cmd_payload_unlocked = 1'b1;
  assign when_Lsu2Plugin_l1698 = (! (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]));
  always @(*) begin
    Lsu2Plugin_logic_special_atomic_loadWhitebox_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
        if(Lsu2Plugin_setup_cacheLoad_rsp_valid) begin
          if(!Lsu2Plugin_setup_cacheLoad_rsp_payload_redo) begin
            if(!Lsu2Plugin_setup_cacheLoad_rsp_payload_fault) begin
              Lsu2Plugin_logic_special_atomic_loadWhitebox_valid = 1'b1;
            end
          end
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_special_atomic_loadWhitebox_readData = Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated[31 : 0];
  always @(*) begin
    Lsu2Plugin_logic_special_atomic_storeWhitebox_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
        Lsu2Plugin_logic_special_atomic_storeWhitebox_valid = 1'b1;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_special_atomic_storeWhitebox_isSc = Lsu2Plugin_logic_special_storeSc;
  assign Lsu2Plugin_logic_special_atomic_storeWhitebox_scPassed = Lsu2Plugin_logic_special_atomic_gotReservation;
  assign FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l1838 = (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]);
  always @(*) begin
    Lsu2Plugin_logic_lqFlush = 1'b0;
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lqFlush = 1'b1;
    end
  end

  assign when_Lsu2Plugin_l1913 = (! Lsu2Plugin_logic_sq_regs_0_commitedNext);
  assign when_Lsu2Plugin_l1913_1 = (! Lsu2Plugin_logic_sq_regs_1_commitedNext);
  assign when_Lsu2Plugin_l1913_2 = (! Lsu2Plugin_logic_sq_regs_2_commitedNext);
  assign when_Lsu2Plugin_l1913_3 = (! Lsu2Plugin_logic_sq_regs_3_commitedNext);
  assign when_Lsu2Plugin_l1913_4 = (! Lsu2Plugin_logic_sq_regs_4_commitedNext);
  assign when_Lsu2Plugin_l1913_5 = (! Lsu2Plugin_logic_sq_regs_5_commitedNext);
  assign when_Lsu2Plugin_l1913_6 = (! Lsu2Plugin_logic_sq_regs_6_commitedNext);
  assign when_Lsu2Plugin_l1913_7 = (! Lsu2Plugin_logic_sq_regs_7_commitedNext);
  assign sqAlloc_0_valid = ((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && FrontendPlugin_dispatch_SQ_ALLOC_0);
  assign sqAlloc_0_id = FrontendPlugin_dispatch_SQ_ID_0;
  assign sqFree_valid = Lsu2Plugin_logic_sq_ptr_onFree_valid;
  assign sqFree_payload = Lsu2Plugin_logic_sq_ptr_onFree_payload;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken = BranchContextPlugin_logic_mem_earlyBranch_spinal_port1;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken[0];
  assign EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken[32 : 1];
  assign EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET = (EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc != EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE);
  assign EU0_BranchPlugin_setup_intFormatPort_payload = _zz_EU0_BranchPlugin_setup_intFormatPort_payload;
  assign EU0_BranchPlugin_logic_branch_badEarlyTaken = (EU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken != EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED = (EU0_BranchPlugin_logic_branch_badEarlyTaken || (EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND && EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET));
  assign EU0_BranchPlugin_setup_reschedule_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  assign EU0_BranchPlugin_setup_reschedule_payload_pcTarget = EU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  assign EU0_BranchPlugin_setup_reschedule_payload_reason = {3'd0, _zz_EU0_BranchPlugin_setup_reschedule_payload_reason};
  assign EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED = ((EU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET[1 : 0] != 2'b00) && EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_isFireing = (EU0_ExecutionUnitBase_pipeline_execute_1_valid && EU0_ExecutionUnitBase_pipeline_execute_1_ready);
  assign EU0_BranchPlugin_setup_reschedule_valid = ((EU0_ExecutionUnitBase_pipeline_execute_1_isFireing && EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL) && (EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED || EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED));
  assign EU0_BranchPlugin_setup_reschedule_payload_trap = EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  assign EU0_BranchPlugin_setup_reschedule_payload_skipCommit = EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  assign EU0_BranchPlugin_setup_reschedule_payload_cause = 4'b0000;
  assign EU0_BranchPlugin_setup_reschedule_payload_tval = EU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  assign EU0_BranchPlugin_logic_branch_finalBranch_valid = (EU0_ExecutionUnitBase_pipeline_execute_1_valid && EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL);
  assign EU0_BranchPlugin_logic_branch_finalBranch_payload_address = EU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID;
  assign EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice = (EU0_ExecutionUnitBase_pipeline_execute_1_PC + _zz_EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice);
  assign EU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget = EU0_ExecutionUnitBase_pipeline_execute_1_PC_TRUE;
  assign EU0_BranchPlugin_logic_branch_finalBranch_payload_data_taken = EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  assign MmuPlugin_logic_satpModeWrite = EU0_CsrAccessPlugin_setup_onWriteBits[31 : 31];
  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_refillOngoing = 1'b0;
    if(MmuPlugin_logic_refill_busy) begin
      if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask) begin
        FetchCachePlugin_setup_translationStorage_logic_refillOngoing = 1'b1;
      end
    end
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask = 4'b0000;
    if(when_MmuPlugin_l522) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask = 4'b1111;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask = ((|_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask) ? _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask_1 : 4'b0000);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address = 2'bxx;
    if(when_MmuPlugin_l522) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter[1:0];
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[13 : 12];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(when_MmuPlugin_l522) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_0) || (! MmuPlugin_logic_refill_load_flags_A));
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault = ((! FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault) && 1'b0);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress = 18'bxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 14];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value == 2'b11);
  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflow = (FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc && FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext = (FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value + _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext);
    if(FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willClear) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext = 2'b00;
    end
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask = 2'b00;
    if(when_MmuPlugin_l522) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask = 2'b11;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask = ((|_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask) ? _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask : 2'b00);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address = 2'bxx;
    if(when_MmuPlugin_l522) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter[1:0];
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[23 : 22];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(when_MmuPlugin_l522) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_1) || (! MmuPlugin_logic_refill_load_flags_A));
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault = ((! FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault) && 1'b0);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress = 8'bxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 24];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress = 10'bxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd22);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc = (FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value == 1'b1);
  assign FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflow = (FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc && FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement);
  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_valueNext = (FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value + FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement);
    if(FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willClear) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_valueNext = 1'b0;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_refillOngoing = 1'b0;
    if(MmuPlugin_logic_refill_busy) begin
      if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask) begin
        Lsu2Plugin_setup_translationStorage_logic_refillOngoing = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask = 4'b0000;
    if(when_MmuPlugin_l522) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask = 4'b1111;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask = ((|_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask) ? _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask_1 : 4'b0000);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address = 2'bxx;
    if(when_MmuPlugin_l522) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter[1:0];
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[13 : 12];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(when_MmuPlugin_l522) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_0) || (! MmuPlugin_logic_refill_load_flags_A));
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault = ((! Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault) && 1'b0);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress = 18'bxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 14];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value == 2'b11);
  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflow = (Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc && Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext = (Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value + _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext);
    if(Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willClear) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext = 2'b00;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask = 2'b00;
    if(when_MmuPlugin_l522) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask = 2'b11;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask = ((|_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask) ? _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask : 2'b00);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address = 2'bxx;
    if(when_MmuPlugin_l522) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter[1:0];
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[23 : 22];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(when_MmuPlugin_l522) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_1) || (! MmuPlugin_logic_refill_load_flags_A));
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault = ((! Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault) && 1'b0);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress = 8'bxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 24];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress = 10'bxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd22);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l499) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc = (Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value == 1'b1);
  assign Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflow = (Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc && Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement);
  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_valueNext = (Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value + Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement);
    if(Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willClear) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_valueNext = 1'b0;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL = Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL_overloaded = ((Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL && (! Lsu2Plugin_setup_translationStorage_logic_refillOngoing)) && Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg);
  assign when_MmuPlugin_l278 = (Lsu2Plugin_logic_sharedPip_stages_0_isRemoved || (! (Lsu2Plugin_logic_sharedPip_stages_0_valid && (! Lsu2Plugin_logic_sharedPip_stages_0_ready))));
  assign Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded = ((Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL && (! Lsu2Plugin_setup_translationStorage_logic_refillOngoing)) && Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg);
  assign when_MmuPlugin_l278_1 = (Lsu2Plugin_logic_sharedPip_stages_1_isRemoved || (! (Lsu2Plugin_logic_sharedPip_stages_1_valid && (! Lsu2Plugin_logic_sharedPip_stages_1_ready))));
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress = Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[13 : 12];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[20 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[40 : 21];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[41];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[42];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[43];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[44];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID[0] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 14]);
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID[1] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 14]);
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID[2] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 14]);
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID[3] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 14]);
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS[0] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID[0] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_valid);
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS[1] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID[1] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_valid);
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS[2] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID[2] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_valid);
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS[3] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID[3] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_valid);
  end

  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[20 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[40 : 21];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[41];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[42];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[43];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[44];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[20 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[40 : 21];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[41];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[42];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[43];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[44];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[20 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[40 : 21];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[41];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[42];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[43];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[44];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_read_1_readAddress = Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[23 : 22];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid = Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[10 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[20 : 11];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[21];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[22];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[23];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[24];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_HITS_PRE_VALID[0] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 24]);
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_HITS_PRE_VALID[1] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 24]);
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS[0] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS_PRE_VALID[0] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_valid);
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS[1] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS_PRE_VALID[1] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_valid);
  end

  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid = Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_spinal_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[10 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[20 : 11];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[21];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[22];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[23];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[24];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS,Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS};
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hit = (|Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits);
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits;
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[1];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[2];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[3];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_4 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[4];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_5 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[5];
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[0] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[1] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[2] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_1));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[3] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_2));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[4] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_4 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_3));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[5] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_5 && (! (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_4 || Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_3)));
  end

  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_1 = (|{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0});
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_2 = (|{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0}});
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_3 = (|{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0}}});
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[0];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[1];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[2];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[3];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[4];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[5];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_6[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated : _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_2) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_3 : _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_5)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_6 : _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_8) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_9 : _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_11))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_12 : 32'h00000000) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_13 : 32'h00000000)));
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault[0];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup = (MmuPlugin_logic_satp_mode == 1'b1);
    if(when_MmuPlugin_l315) begin
      Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
    if(when_MmuPlugin_l316) begin
      if(when_MmuPlugin_l318) begin
        Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
      end
    end
  end

  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_needRefill = ((Lsu2Plugin_logic_sharedPip_stages_1_valid && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hit)) && Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup);
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_askRefill = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_needRefill && Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded);
  assign when_MmuPlugin_l315 = ((! MmuPlugin_logic_status_mprv) && (PrivilegedPlugin_setup_privilege == 2'b11));
  assign when_MmuPlugin_l316 = (PrivilegedPlugin_setup_privilege == 2'b11);
  assign when_MmuPlugin_l318 = ((! MmuPlugin_logic_status_mprv) || (PrivilegedPlugin_logic_machine_mstatus_mpp == 2'b11));
  assign EU0_CsrAccessPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_wantStart = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
        EU0_CsrAccessPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign EU0_CsrAccessPlugin_logic_fsm_wantKill = 1'b0;
  assign CsrRamPlugin_logic_flush_done = CsrRamPlugin_logic_flush_counter[3];
  assign CsrRamPlugin_setup_initPort_valid = (! CsrRamPlugin_logic_flush_done);
  assign CsrRamPlugin_setup_initPort_address = CsrRamPlugin_logic_flush_counter[2:0];
  assign CsrRamPlugin_setup_initPort_data = 32'h00000000;
  assign when_CsrRamPlugin_l61 = ((! CsrRamPlugin_logic_flush_done) && CsrRamPlugin_setup_initPort_ready);
  assign CsrRamPlugin_logic_writeLogic_hits = {CsrRamPlugin_setup_initPort_valid,{PrivilegedPlugin_setup_ramWrite_valid,EU0_CsrAccessPlugin_logic_ramWritePort_valid}};
  assign CsrRamPlugin_logic_writeLogic_hit = (|CsrRamPlugin_logic_writeLogic_hits);
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_input = CsrRamPlugin_logic_writeLogic_hits;
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_writeLogic_oh = CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  assign _zz_PrivilegedPlugin_setup_ramWrite_ready = CsrRamPlugin_logic_writeLogic_oh[1];
  assign _zz_CsrRamPlugin_setup_initPort_ready = CsrRamPlugin_logic_writeLogic_oh[2];
  assign CsrRamPlugin_logic_writeLogic_sel = {_zz_CsrRamPlugin_setup_initPort_ready,_zz_PrivilegedPlugin_setup_ramWrite_ready};
  assign CsrRamPlugin_logic_writeLogic_port_valid = CsrRamPlugin_logic_writeLogic_hit;
  assign CsrRamPlugin_logic_writeLogic_port_payload_address = _zz_CsrRamPlugin_logic_writeLogic_port_payload_address;
  assign CsrRamPlugin_logic_writeLogic_port_payload_data = _zz_CsrRamPlugin_logic_writeLogic_port_payload_data;
  assign EU0_CsrAccessPlugin_logic_ramWritePort_ready = CsrRamPlugin_logic_writeLogic_oh[0];
  assign PrivilegedPlugin_setup_ramWrite_ready = _zz_PrivilegedPlugin_setup_ramWrite_ready;
  assign CsrRamPlugin_setup_initPort_ready = _zz_CsrRamPlugin_setup_initPort_ready;
  assign CsrRamPlugin_logic_readLogic_hits = {PrivilegedPlugin_setup_ramRead_valid,EU0_CsrAccessPlugin_logic_ramReadPort_valid};
  assign CsrRamPlugin_logic_readLogic_hit = (|CsrRamPlugin_logic_readLogic_hits);
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_input = CsrRamPlugin_logic_readLogic_hits;
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_readLogic_oh = CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  assign _zz_PrivilegedPlugin_setup_ramRead_ready = CsrRamPlugin_logic_readLogic_oh[1];
  assign CsrRamPlugin_logic_readLogic_sel = _zz_PrivilegedPlugin_setup_ramRead_ready;
  assign CsrRamPlugin_logic_readLogic_port_data = CsrRamPlugin_logic_mem_spinal_port1;
  assign CsrRamPlugin_logic_readLogic_port_address = _zz_CsrRamPlugin_logic_readLogic_port_address;
  assign EU0_CsrAccessPlugin_logic_ramReadPort_ready = CsrRamPlugin_logic_readLogic_oh[0];
  assign PrivilegedPlugin_setup_ramRead_ready = _zz_PrivilegedPlugin_setup_ramRead_ready;
  assign EU0_CsrAccessPlugin_logic_ramReadPort_data = CsrRamPlugin_logic_readLogic_port_data;
  assign PrivilegedPlugin_setup_ramRead_data = CsrRamPlugin_logic_readLogic_port_data;
  always @(*) begin
    PrivilegedPlugin_setup_ramWrite_valid = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_ramWrite_address = 3'bxxx;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_address = _zz_PrivilegedPlugin_setup_ramWrite_address;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_address = _zz_PrivilegedPlugin_setup_ramWrite_address_1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_ramWrite_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_data = _zz_PrivilegedPlugin_setup_ramWrite_data;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_data = _zz_PrivilegedPlugin_setup_ramWrite_data_1;
        if(PrivilegedPlugin_logic_decoderInterrupt_raised) begin
          PrivilegedPlugin_setup_ramWrite_data = 32'h00000000;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_ramRead_valid = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        PrivilegedPlugin_setup_ramRead_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        PrivilegedPlugin_setup_ramRead_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_ramRead_address = 3'bxxx;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        PrivilegedPlugin_setup_ramRead_address = _zz_PrivilegedPlugin_setup_ramRead_address;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        PrivilegedPlugin_setup_ramRead_address = _zz_PrivilegedPlugin_setup_ramRead_address_1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_logic_interrupt_valid = 1'b0;
    if(when_PrivilegedPlugin_l638_1) begin
      if(when_PrivilegedPlugin_l644) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l644_1) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l644_2) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
    end
    if(when_PrivilegedPlugin_l638) begin
      if(when_PrivilegedPlugin_l644_3) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l644_4) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l644_5) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l644_6) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l644_7) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l644_8) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_interrupt_code = 4'bxxxx;
    if(when_PrivilegedPlugin_l638_1) begin
      if(when_PrivilegedPlugin_l644) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0001;
      end
      if(when_PrivilegedPlugin_l644_1) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0101;
      end
      if(when_PrivilegedPlugin_l644_2) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b1001;
      end
    end
    if(when_PrivilegedPlugin_l638) begin
      if(when_PrivilegedPlugin_l644_3) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0111;
      end
      if(when_PrivilegedPlugin_l644_4) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0011;
      end
      if(when_PrivilegedPlugin_l644_5) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b1011;
      end
      if(when_PrivilegedPlugin_l644_6) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0001;
      end
      if(when_PrivilegedPlugin_l644_7) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0101;
      end
      if(when_PrivilegedPlugin_l644_8) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b1001;
      end
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'bxx;
    if(when_PrivilegedPlugin_l638_1) begin
      if(when_PrivilegedPlugin_l644) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b01;
      end
      if(when_PrivilegedPlugin_l644_1) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b01;
      end
      if(when_PrivilegedPlugin_l644_2) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b01;
      end
    end
    if(when_PrivilegedPlugin_l638) begin
      if(when_PrivilegedPlugin_l644_3) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l644_4) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l644_5) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l644_6) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l644_7) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l644_8) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
    end
  end

  assign when_PrivilegedPlugin_l638 = (PrivilegedPlugin_logic_machine_mstatus_mie || (! PrivilegedPlugin_setup_withMachinePrivilege));
  assign when_PrivilegedPlugin_l638_1 = ((PrivilegedPlugin_logic_supervisor_sstatus_sie && (! PrivilegedPlugin_setup_withMachinePrivilege)) || (! PrivilegedPlugin_setup_withSupervisorPrivilege));
  assign when_PrivilegedPlugin_l644 = ((_zz_when_PrivilegedPlugin_l644 && (1'b1 && PrivilegedPlugin_logic_machine_mideleg_ss)) && (! 1'b0));
  assign when_PrivilegedPlugin_l644_1 = ((_zz_when_PrivilegedPlugin_l644_1 && (1'b1 && PrivilegedPlugin_logic_machine_mideleg_st)) && (! 1'b0));
  assign when_PrivilegedPlugin_l644_2 = ((_zz_when_PrivilegedPlugin_l644_2 && (1'b1 && PrivilegedPlugin_logic_machine_mideleg_se)) && (! 1'b0));
  assign when_PrivilegedPlugin_l644_3 = (((PrivilegedPlugin_logic_machine_mip_mtip && PrivilegedPlugin_logic_machine_mie_mtie) && 1'b1) && (! 1'b0));
  assign when_PrivilegedPlugin_l644_4 = (((PrivilegedPlugin_logic_machine_mip_msip && PrivilegedPlugin_logic_machine_mie_msie) && 1'b1) && (! 1'b0));
  assign when_PrivilegedPlugin_l644_5 = (((PrivilegedPlugin_logic_machine_mip_meip && PrivilegedPlugin_logic_machine_mie_meie) && 1'b1) && (! 1'b0));
  assign when_PrivilegedPlugin_l644_6 = ((_zz_when_PrivilegedPlugin_l644 && 1'b1) && (! (|PrivilegedPlugin_logic_machine_mideleg_ss)));
  assign when_PrivilegedPlugin_l644_7 = ((_zz_when_PrivilegedPlugin_l644_1 && 1'b1) && (! (|PrivilegedPlugin_logic_machine_mideleg_st)));
  assign when_PrivilegedPlugin_l644_8 = ((_zz_when_PrivilegedPlugin_l644_2 && 1'b1) && (! (|PrivilegedPlugin_logic_machine_mideleg_se)));
  assign PrivilegedPlugin_logic_decoderInterrupt_doIt = PrivilegedPlugin_logic_decoderInterrupt_counter[2];
  assign when_PrivilegedPlugin_l675 = (((! PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt) || (! DecoderPlugin_setup_trapReady)) || PrivilegedPlugin_logic_decoderInterrupt_raised);
  assign when_PrivilegedPlugin_l679 = (PrivilegedPlugin_logic_decoderInterrupt_doIt && (! PrivilegedPlugin_logic_decoderInterrupt_raised));
  assign PrivilegedPlugin_logic_decoderInterrupt_buffer_sample = (PrivilegedPlugin_logic_interrupt_valid && (! PrivilegedPlugin_logic_decoderInterrupt_raised));
  always @(*) begin
    PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b11;
    case(PrivilegedPlugin_logic_exception_code)
      4'b0000 : begin
        if(when_PrivilegedPlugin_l709) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b0011 : begin
        if(when_PrivilegedPlugin_l709_1) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1000 : begin
        if(when_PrivilegedPlugin_l709_2) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1001 : begin
        if(when_PrivilegedPlugin_l709_3) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1100 : begin
        if(when_PrivilegedPlugin_l709_4) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1101 : begin
        if(when_PrivilegedPlugin_l709_5) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1111 : begin
        if(when_PrivilegedPlugin_l709_6) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_logic_exception_code = PrivilegedPlugin_logic_reschedule_payload_cause;
    if(when_PrivilegedPlugin_l696) begin
      PrivilegedPlugin_logic_exception_code[1 : 0] = PrivilegedPlugin_setup_privilege;
    end
  end

  assign when_PrivilegedPlugin_l696 = (PrivilegedPlugin_logic_reschedule_payload_cause == 4'b1011);
  assign when_PrivilegedPlugin_l709 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_iam) && (! 1'b0));
  assign when_PrivilegedPlugin_l709_1 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_bp) && (! 1'b0));
  assign when_PrivilegedPlugin_l709_2 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_eu) && (! 1'b0));
  assign when_PrivilegedPlugin_l709_3 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_es) && (! 1'b0));
  assign when_PrivilegedPlugin_l709_4 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_ipf) && (! 1'b0));
  assign when_PrivilegedPlugin_l709_5 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_lpf) && (! 1'b0));
  assign when_PrivilegedPlugin_l709_6 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_spf) && (! 1'b0));
  assign PrivilegedPlugin_logic_exception_targetPrivilege = ((PrivilegedPlugin_setup_privilege < PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped) ? PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped : PrivilegedPlugin_setup_privilege);
  assign PrivilegedPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    PrivilegedPlugin_logic_fsm_wantStart = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
        PrivilegedPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign PrivilegedPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    PrivilegedPlugin_logic_fsm_trap_fire = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_logic_fsm_trap_fire = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_logic_fsm_xret_sourcePrivilege = PrivilegedPlugin_logic_reschedule_payload_tval[1 : 0];
  always @(*) begin
    PrivilegedPlugin_logic_fsm_xret_targetPrivilege = PrivilegedPlugin_logic_machine_mstatus_mpp;
    case(PrivilegedPlugin_logic_fsm_xret_sourcePrivilege)
      2'b01 : begin
        PrivilegedPlugin_logic_fsm_xret_targetPrivilege = {1'b0,PrivilegedPlugin_logic_supervisor_sstatus_spp};
      end
      default : begin
      end
    endcase
  end

  assign FetchPlugin_stages_0_haltRequest_PrivilegedPlugin_l975 = ((! (PrivilegedPlugin_logic_fsm_stateReg == PrivilegedPlugin_logic_fsm_enumDef_IDLE)) || (CommitPlugin_logic_reschedule_valid && CommitPlugin_logic_reschedule_trap));
  assign trap_fire = PrivilegedPlugin_logic_fsm_trap_fire;
  assign trap_code = PrivilegedPlugin_logic_fsm_trap_code;
  assign trap_interrupt = PrivilegedPlugin_logic_fsm_trap_interrupt;
  assign trap_tval = PrivilegedPlugin_logic_reschedule_payload_tval;
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_immZero = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[19 : 15] == 5'h00);
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_srcZero = (EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_IMM ? EU0_CsrAccessPlugin_logic_fsm_startLogic_immZero : (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[19 : 15] == 5'h00));
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_csrWrite = (! (EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK && EU0_CsrAccessPlugin_logic_fsm_startLogic_srcZero));
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_csrRead = (! ((! EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK) && (! EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD)));
  assign COMB_CSR_773 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h305);
  assign COMB_CSR_835 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h343);
  assign COMB_CSR_833 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h341);
  assign COMB_CSR_832 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h340);
  assign COMB_CSR_3857 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hf11);
  assign COMB_CSR_3858 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hf12);
  assign COMB_CSR_3859 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hf13);
  assign COMB_CSR_3860 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hf14);
  assign COMB_CSR_769 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h301);
  assign COMB_CSR_834 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h342);
  assign COMB_CSR_768 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h300);
  assign COMB_CSR_836 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h344);
  assign COMB_CSR_772 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h304);
  assign COMB_CSR_770 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h302);
  assign COMB_CSR_771 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h303);
  assign COMB_CSR_261 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h105);
  assign COMB_CSR_323 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h143);
  assign COMB_CSR_321 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h141);
  assign COMB_CSR_320 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h140);
  assign COMB_CSR_322 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h142);
  assign COMB_CSR_256 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h100);
  assign COMB_CSR_260 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h104);
  assign COMB_CSR_324 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h144);
  assign COMB_CSR_384 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h180);
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented = (|{COMB_CSR_384,{COMB_CSR_324,{COMB_CSR_260,{COMB_CSR_256,{COMB_CSR_322,{COMB_CSR_320,{COMB_CSR_321,{COMB_CSR_323,{COMB_CSR_261,{COMB_CSR_771,{_zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented,_zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_1}}}}}}}}}}});
  assign EU0_CsrAccessPlugin_setup_onDecodeWrite = EU0_CsrAccessPlugin_logic_fsm_startLogic_csrWrite;
  assign EU0_CsrAccessPlugin_setup_onDecodeRead = EU0_CsrAccessPlugin_logic_fsm_startLogic_csrRead;
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_trap = ((! EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented) || EU0_CsrAccessPlugin_setup_onDecodeTrap);
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_write = ((EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL && (! EU0_CsrAccessPlugin_logic_fsm_startLogic_trap)) && EU0_CsrAccessPlugin_logic_fsm_startLogic_csrWrite);
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_read = ((EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL && (! EU0_CsrAccessPlugin_logic_fsm_startLogic_trap)) && EU0_CsrAccessPlugin_logic_fsm_startLogic_csrRead);
  assign EU0_CsrAccessPlugin_setup_onDecodeAddress = _zz_EU0_CsrAccessPlugin_setup_onDecodeAddress[31 : 20];
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_onDecodeDo = (EU0_ExecutionUnitBase_pipeline_execute_0_valid && EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL);
  assign when_CsrAccessPlugin_l183 = (EU0_CsrAccessPlugin_logic_fsm_startLogic_onDecodeDo && COMB_CSR_384);
  assign when_MmuPlugin_l218 = (PrivilegedPlugin_logic_machine_mstatus_tvm && (PrivilegedPlugin_setup_privilege == 2'b01));
  assign EU0_CsrAccessPlugin_setup_onReadAddress = _zz_EU0_CsrAccessPlugin_setup_onReadAddress[31 : 20];
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = EU0_CsrAccessPlugin_logic_fsm_regs_read;
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        if(when_CsrAccessPlugin_l285) begin
          EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = EU0_CsrAccessPlugin_logic_fsm_regs_read;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign EU0_CsrAccessPlugin_setup_onReadMovingOff = ((! EU0_CsrAccessPlugin_setup_onReadHalt) || EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed);
  assign _zz_259 = zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue(1'b0);
  always @(*) _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue = _zz_259;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1[31 : 0] = 32'h40141101;
  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2[31 : 31] = PrivilegedPlugin_logic_machine_cause_interrupt;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2[3 : 0] = PrivilegedPlugin_logic_machine_cause_code;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[12 : 11] = PrivilegedPlugin_logic_machine_mstatus_mpp;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[7 : 7] = PrivilegedPlugin_logic_machine_mstatus_mpie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[3 : 3] = PrivilegedPlugin_logic_machine_mstatus_mie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[31 : 31] = PrivilegedPlugin_logic_machine_mstatus_sd;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[22 : 22] = PrivilegedPlugin_logic_machine_mstatus_tsr;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[21 : 21] = PrivilegedPlugin_logic_machine_mstatus_tw;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[20 : 20] = PrivilegedPlugin_logic_machine_mstatus_tvm;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[14 : 13] = PrivilegedPlugin_logic_machine_mstatus_fs;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[8 : 8] = PrivilegedPlugin_logic_supervisor_sstatus_spp;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[5 : 5] = PrivilegedPlugin_logic_supervisor_sstatus_spie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[1 : 1] = PrivilegedPlugin_logic_supervisor_sstatus_sie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[19 : 19] = MmuPlugin_logic_status_mxr;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[18 : 18] = MmuPlugin_logic_status_sum;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[17 : 17] = MmuPlugin_logic_status_mprv;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[11 : 11] = PrivilegedPlugin_logic_machine_mip_meip;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[7 : 7] = PrivilegedPlugin_logic_machine_mip_mtip;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[3 : 3] = PrivilegedPlugin_logic_machine_mip_msip;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[9 : 9] = PrivilegedPlugin_logic_supervisor_sip_seipOr;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[5 : 5] = PrivilegedPlugin_logic_supervisor_sip_stip;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[1 : 1] = PrivilegedPlugin_logic_supervisor_sip_ssip;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[11 : 11] = PrivilegedPlugin_logic_machine_mie_meie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[7 : 7] = PrivilegedPlugin_logic_machine_mie_mtie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[3 : 3] = PrivilegedPlugin_logic_machine_mie_msie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[9 : 9] = PrivilegedPlugin_logic_supervisor_sie_seie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[5 : 5] = PrivilegedPlugin_logic_supervisor_sie_stie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[1 : 1] = PrivilegedPlugin_logic_supervisor_sie_ssie;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[0 : 0] = PrivilegedPlugin_logic_machine_medeleg_iam;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[3 : 3] = PrivilegedPlugin_logic_machine_medeleg_bp;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[8 : 8] = PrivilegedPlugin_logic_machine_medeleg_eu;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[9 : 9] = PrivilegedPlugin_logic_machine_medeleg_es;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[12 : 12] = PrivilegedPlugin_logic_machine_medeleg_ipf;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[13 : 13] = PrivilegedPlugin_logic_machine_medeleg_lpf;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[15 : 15] = PrivilegedPlugin_logic_machine_medeleg_spf;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7[9 : 9] = PrivilegedPlugin_logic_machine_mideleg_se;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7[5 : 5] = PrivilegedPlugin_logic_machine_mideleg_st;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7[1 : 1] = PrivilegedPlugin_logic_machine_mideleg_ss;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8[31 : 31] = PrivilegedPlugin_logic_supervisor_cause_interrupt;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8[3 : 0] = PrivilegedPlugin_logic_supervisor_cause_code;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[8 : 8] = PrivilegedPlugin_logic_supervisor_sstatus_spp;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[5 : 5] = PrivilegedPlugin_logic_supervisor_sstatus_spie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[1 : 1] = PrivilegedPlugin_logic_supervisor_sstatus_sie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[14 : 13] = PrivilegedPlugin_logic_machine_mstatus_fs;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[31 : 31] = PrivilegedPlugin_logic_machine_mstatus_sd;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[19 : 19] = MmuPlugin_logic_status_mxr;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[18 : 18] = MmuPlugin_logic_status_sum;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10[9 : 9] = (PrivilegedPlugin_logic_supervisor_sie_seie && PrivilegedPlugin_logic_machine_mideleg_se);
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10[5 : 5] = (PrivilegedPlugin_logic_supervisor_sie_stie && PrivilegedPlugin_logic_machine_mideleg_st);
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10[1 : 1] = (PrivilegedPlugin_logic_supervisor_sie_ssie && PrivilegedPlugin_logic_machine_mideleg_ss);
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11[9 : 9] = (PrivilegedPlugin_logic_supervisor_sip_seipOr && PrivilegedPlugin_logic_machine_mideleg_se);
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11[5 : 5] = (PrivilegedPlugin_logic_supervisor_sip_stip && PrivilegedPlugin_logic_machine_mideleg_st);
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11[1 : 1] = (PrivilegedPlugin_logic_supervisor_sip_ssip && PrivilegedPlugin_logic_machine_mideleg_ss);
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12[31 : 31] = MmuPlugin_logic_satp_mode;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12[19 : 0] = MmuPlugin_logic_satp_ppn;
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue = (((((REG_CSR_3857 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14) | (REG_CSR_3858 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15)) | ((REG_CSR_3859 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17) | (REG_CSR_3860 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19))) | (((REG_CSR_769 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20) | (REG_CSR_834 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21)) | ((REG_CSR_768 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22) | (REG_CSR_836 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23)))) | ((((REG_CSR_772 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24) | (REG_CSR_770 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25)) | ((REG_CSR_771 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26) | (REG_CSR_322 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27))) | (((REG_CSR_256 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28) | (REG_CSR_260 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29)) | ((REG_CSR_324 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30) | (REG_CSR_384 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31)))));
    if(EU0_CsrAccessPlugin_logic_fsm_regs_ramSel) begin
      EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue = EU0_CsrAccessPlugin_logic_ramReadPort_data;
    end
  end

  assign EU0_CsrAccessPlugin_logic_ramReadPort_valid = (EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && EU0_CsrAccessPlugin_logic_fsm_regs_ramSel);
  assign EU0_CsrAccessPlugin_logic_ramReadPort_address = EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress;
  assign when_CsrAccessPlugin_l272 = (EU0_CsrAccessPlugin_logic_ramReadPort_valid && (! EU0_CsrAccessPlugin_logic_ramReadPort_ready));
  always @(*) begin
    EU0_CsrAccessPlugin_setup_onReadToWriteBits = EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
    if(when_CsrAccessPlugin_l278) begin
      EU0_CsrAccessPlugin_setup_onReadToWriteBits[9 : 9] = PrivilegedPlugin_logic_supervisor_sip_seipSoft;
    end
  end

  assign when_CsrAccessPlugin_l278 = (EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_836);
  assign EU0_CsrAccessPlugin_setup_onWriteMovingOff = ((! EU0_CsrAccessPlugin_setup_onWriteHalt) || EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed);
  assign EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = (EU0_CsrAccessPlugin_logic_fsm_regs_doImm ? _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask : EU0_CsrAccessPlugin_logic_fsm_regs_rs1);
  assign EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_masked = (EU0_CsrAccessPlugin_logic_fsm_regs_doClear ? (EU0_CsrAccessPlugin_logic_fsm_regs_aluInput & (~ EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask)) : (EU0_CsrAccessPlugin_logic_fsm_regs_aluInput | EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask));
  assign EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_result = (EU0_CsrAccessPlugin_logic_fsm_regs_doMask ? EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_masked : EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask);
  always @(*) begin
    EU0_CsrAccessPlugin_setup_onWriteBits = EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(when_CsrAccessPlugin_l327) begin
      EU0_CsrAccessPlugin_setup_onWriteBits[1 : 0] = 2'b00;
    end
    if(when_CsrAccessPlugin_l327_1) begin
      EU0_CsrAccessPlugin_setup_onWriteBits[1 : 0] = 2'b00;
    end
  end

  assign EU0_CsrAccessPlugin_setup_onWriteAddress = _zz_EU0_CsrAccessPlugin_setup_onWriteAddress[31 : 20];
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = EU0_CsrAccessPlugin_logic_fsm_regs_write;
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        if(when_CsrAccessPlugin_l311) begin
          EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = EU0_CsrAccessPlugin_logic_fsm_regs_write;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign when_CsrAccessPlugin_l327 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_833);
  assign when_CsrAccessPlugin_l328 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_834);
  assign when_CsrAccessPlugin_l328_1 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_768);
  assign when_CsrAccessPlugin_l328_2 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_836);
  assign when_CsrAccessPlugin_l328_3 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_772);
  assign when_CsrAccessPlugin_l328_4 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_770);
  assign when_CsrAccessPlugin_l328_5 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_771);
  assign when_CsrAccessPlugin_l327_1 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_321);
  assign when_CsrAccessPlugin_l328_6 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_322);
  assign when_CsrAccessPlugin_l328_7 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_256);
  assign when_CsrAccessPlugin_l328_8 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_260);
  assign when_CsrAccessPlugin_l328_9 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_324);
  assign when_CsrAccessPlugin_l333 = ((|((MmuPlugin_logic_satpModeWrite != 1'b0) && (MmuPlugin_logic_satpModeWrite != 1'b1))) == 1'b0);
  assign when_CsrAccessPlugin_l328_10 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_384);
  assign when_CsrAccessPlugin_l338 = (EU0_CsrAccessPlugin_logic_ramWritePort_valid && EU0_CsrAccessPlugin_logic_ramWritePort_ready);
  assign EU0_CsrAccessPlugin_logic_ramWritePort_valid = ((EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && EU0_CsrAccessPlugin_logic_fsm_regs_ramSel) && (! EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired));
  assign EU0_CsrAccessPlugin_logic_ramWritePort_address = EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress;
  assign EU0_CsrAccessPlugin_logic_ramWritePort_data = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign when_CsrAccessPlugin_l342 = (EU0_CsrAccessPlugin_logic_ramWritePort_valid && (! EU0_CsrAccessPlugin_logic_ramWritePort_ready));
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_isDone = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
        EU0_CsrAccessPlugin_logic_fsm_isDone = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_isCompletionReady = 1'b0;
    if(EU0_ExecutionUnitBase_pipeline_execute_2_ready) begin
      EU0_CsrAccessPlugin_logic_fsm_isCompletionReady = 1'b1;
    end
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_stateReg;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
        if(EU0_CsrAccessPlugin_logic_fsm_startLogic_onDecodeDo) begin
          EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_READ;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        if(when_CsrAccessPlugin_l285) begin
          EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        if(when_CsrAccessPlugin_l311) begin
          EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
        if(EU0_CsrAccessPlugin_logic_fsm_isCompletionReady) begin
          EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed) begin
      EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE;
    end
    if(EU0_CsrAccessPlugin_logic_fsm_wantStart) begin
      EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE;
    end
    if(EU0_CsrAccessPlugin_logic_fsm_wantKill) begin
      EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT;
    end
  end

  assign switch_CsrAccessPlugin_l206 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign when_CsrAccessPlugin_l285 = (! EU0_CsrAccessPlugin_setup_onReadHalt);
  assign when_CsrAccessPlugin_l311 = (! EU0_CsrAccessPlugin_setup_onWriteHalt);
  assign EU0_CsrAccessPlugin_setup_intFormatPort_payload = EU0_CsrAccessPlugin_logic_fsm_regs_csrValue;
  assign EU0_CsrAccessPlugin_setup_trap_valid = (((EU0_ExecutionUnitBase_pipeline_execute_2_valid && EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL) && EU0_CsrAccessPlugin_logic_fsm_isDone) && (EU0_CsrAccessPlugin_logic_fsm_regs_trap || EU0_CsrAccessPlugin_logic_fsm_regs_flushPipeline));
  assign EU0_CsrAccessPlugin_setup_trap_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  always @(*) begin
    EU0_CsrAccessPlugin_setup_trap_payload_cause = 4'b0010;
    if(when_CsrAccessPlugin_l378) begin
      EU0_CsrAccessPlugin_setup_trap_payload_cause = 4'b1001;
    end
  end

  assign EU0_CsrAccessPlugin_setup_trap_payload_tval = EU0_CsrAccessPlugin_logic_fsm_regs_microOp;
  assign EU0_CsrAccessPlugin_setup_trap_payload_skipCommit = EU0_CsrAccessPlugin_logic_fsm_regs_trap;
  assign EU0_CsrAccessPlugin_setup_trap_payload_reason = 8'h01;
  assign EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_CsrAccessPlugin_l375 = ((EU0_ExecutionUnitBase_pipeline_execute_2_valid && EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL) && (! EU0_CsrAccessPlugin_logic_fsm_isDone));
  assign when_CsrAccessPlugin_l378 = (! EU0_CsrAccessPlugin_logic_fsm_regs_trap);
  assign EU0_ExecutionUnitBase_pipeline_execute_2_isFireing = (EU0_ExecutionUnitBase_pipeline_execute_2_valid && EU0_ExecutionUnitBase_pipeline_execute_2_ready);
  assign csrAccess_valid = ((EU0_ExecutionUnitBase_pipeline_execute_2_isFireing && EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL) && (! EU0_CsrAccessPlugin_logic_fsm_regs_trap));
  assign csrAccess_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  assign csrAccess_payload_address = _zz_csrAccess_payload_address[31 : 20];
  assign csrAccess_payload_write = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign csrAccess_payload_read = EU0_CsrAccessPlugin_logic_fsm_regs_csrValue;
  assign csrAccess_payload_writeDone = EU0_CsrAccessPlugin_logic_fsm_regs_write;
  assign csrAccess_payload_readDone = EU0_CsrAccessPlugin_logic_fsm_regs_read;
  assign csrAccess_payload_fsDirty = 1'b0;
  assign EnvCallPlugin_setup_reschedule_valid = (EU0_ExecutionUnitBase_pipeline_execute_2_valid && ((((((EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA) || (EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_WFI && (! ((PrivilegedPlugin_setup_privilege == 2'b11) || ((! PrivilegedPlugin_logic_machine_mstatus_tw) && (1'b0 || (PrivilegedPlugin_setup_privilege == 2'b01))))))));
  assign EnvCallPlugin_setup_reschedule_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  always @(*) begin
    EnvCallPlugin_setup_reschedule_payload_tval = (EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK ? EU0_ExecutionUnitBase_pipeline_execute_2_PC : 32'h00000000);
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) begin
      EnvCallPlugin_setup_reschedule_payload_tval[1 : 0] = EnvCallPlugin_logic_xretPriv;
    end
  end

  always @(*) begin
    EnvCallPlugin_setup_reschedule_payload_skipCommit = (EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL);
    if(EnvCallPlugin_logic_trap) begin
      EnvCallPlugin_setup_reschedule_payload_skipCommit = 1'b1;
    end
  end

  always @(*) begin
    EnvCallPlugin_setup_reschedule_payload_reason = 8'h02;
    if(EnvCallPlugin_logic_trap) begin
      EnvCallPlugin_setup_reschedule_payload_reason = 8'h01;
    end
  end

  always @(*) begin
    EnvCallPlugin_setup_reschedule_payload_cause = 4'bxxxx;
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b1000;
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b0011;
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b1011;
    end
    if(when_EnvCallPlugin_l108) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b1001;
    end
    if(EnvCallPlugin_logic_trap) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b0010;
    end
  end

  assign EnvCallPlugin_logic_xretPriv = EU0_ExecutionUnitBase_pipeline_execute_2_Frontend_MICRO_OP[29 : 28];
  always @(*) begin
    EnvCallPlugin_logic_trap = 1'b0;
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) begin
      if(when_EnvCallPlugin_l99) begin
        EnvCallPlugin_logic_trap = 1'b1;
      end
      if(when_EnvCallPlugin_l100) begin
        EnvCallPlugin_logic_trap = 1'b1;
      end
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA) begin
      if(when_EnvCallPlugin_l112) begin
        EnvCallPlugin_logic_trap = 1'b1;
      end
      if(when_EnvCallPlugin_l113) begin
        EnvCallPlugin_logic_trap = 1'b1;
      end
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_WFI) begin
      EnvCallPlugin_logic_trap = 1'b1;
    end
  end

  assign when_EnvCallPlugin_l99 = (PrivilegedPlugin_setup_privilege < EnvCallPlugin_logic_xretPriv);
  assign when_EnvCallPlugin_l100 = ((PrivilegedPlugin_logic_machine_mstatus_tsr && (PrivilegedPlugin_setup_privilege == 2'b01)) && (EnvCallPlugin_logic_xretPriv == 2'b01));
  assign when_EnvCallPlugin_l108 = ((EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA);
  assign when_EnvCallPlugin_l112 = ((PrivilegedPlugin_setup_privilege == 2'b01) && PrivilegedPlugin_logic_machine_mstatus_tvm);
  assign when_EnvCallPlugin_l113 = (PrivilegedPlugin_setup_privilege == 2'b00);
  assign EnvCallPlugin_logic_flushes_wantExit = 1'b0;
  always @(*) begin
    EnvCallPlugin_logic_flushes_wantStart = 1'b0;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
        EnvCallPlugin_logic_flushes_wantStart = 1'b1;
      end
    endcase
  end

  assign EnvCallPlugin_logic_flushes_wantKill = 1'b0;
  assign FetchPlugin_stages_0_haltRequest_EnvCallPlugin_l138 = (! (EnvCallPlugin_logic_flushes_stateReg == EnvCallPlugin_logic_flushes_enumDef_IDLE));
  always @(*) begin
    EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_stateReg;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
        if(EU0_ExecutionUnitBase_pipeline_execute_2_valid) begin
          if(EU0_ExecutionUnitBase_pipeline_execute_2_ready) begin
            if(when_EnvCallPlugin_l148) begin
              EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE;
            end
            if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA) begin
              EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH;
            end
          end
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
        if(CommitPlugin_logic_commit_reschedulePort_valid) begin
          EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
        EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT;
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
        if(FetchCachePlugin_setup_invalidatePort_rsp_valid) begin
          EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH;
        end
        if(MmuPlugin_setup_invalidatePort_rsp_valid) begin
          EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_IDLE;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
        EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU;
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
        if(Lsu2Plugin_setup_flushPort_rsp_valid) begin
          EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(EnvCallPlugin_logic_flushes_wantStart) begin
      EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_IDLE;
    end
    if(EnvCallPlugin_logic_flushes_wantKill) begin
      EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_BOOT;
    end
  end

  assign when_EnvCallPlugin_l148 = (EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA);
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO = ((ioStartAddr <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED) && (Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED <= _zz_FetchPlugin_stages_1_MMU_IO));
  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO = (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hit);
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO = 1'b0;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_EXECUTE = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute && (! (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser && (PrivilegedPlugin_setup_privilege == 2'b01))));
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_EXECUTE = 1'b1;
    end
    if(when_MmuPlugin_l356) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_EXECUTE = 1'b0;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ = 1'b1;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_WRITE = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_WRITE = 1'b1;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT = ((Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException || ((Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser && (PrivilegedPlugin_setup_privilege == 2'b01)) && (! MmuPlugin_logic_status_sum))) || ((! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser) && (PrivilegedPlugin_setup_privilege == 2'b00)));
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT = 1'b0;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT = (1'b0 || (! (1'b1 || Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO)));
    end
  end

  assign when_MmuPlugin_l356 = (! 1'b1);
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_BYPASS_TRANSLATION = (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup);
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_OH = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh;
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_0 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_1 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_2 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_3 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_4 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[21 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_5 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[21 : 0]};
  assign FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL = 1'b1;
  assign FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded = ((FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL && (! FetchCachePlugin_setup_translationStorage_logic_refillOngoing)) && FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg);
  assign when_MmuPlugin_l278_2 = (FetchPlugin_stages_1_isRemoved || (! (FetchPlugin_stages_1_valid && (! FetchPlugin_stages_1_ready))));
  assign FetchCachePlugin_logic_translationPort_logic_read_0_readAddress = FetchPlugin_stages_1_Fetch_FETCH_PC[13 : 12];
  assign _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_spinal_port1;
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[0];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_pageFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[1];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_accessFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[2];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[20 : 3];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[40 : 21];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowRead = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[41];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowWrite = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[42];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowExecute = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[43];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowUser = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[44];
  always @(*) begin
    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[0] = (FetchPlugin_stages_1_MMU_L0_ENTRIES_0_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 14]);
    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[1] = (FetchPlugin_stages_1_MMU_L0_ENTRIES_1_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 14]);
    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[2] = (FetchPlugin_stages_1_MMU_L0_ENTRIES_2_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 14]);
    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[3] = (FetchPlugin_stages_1_MMU_L0_ENTRIES_3_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 14]);
  end

  always @(*) begin
    FetchPlugin_stages_1_MMU_L0_HITS[0] = (FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[0] && FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid);
    FetchPlugin_stages_1_MMU_L0_HITS[1] = (FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[1] && FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid);
    FetchPlugin_stages_1_MMU_L0_HITS[2] = (FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[2] && FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid);
    FetchPlugin_stages_1_MMU_L0_HITS[3] = (FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[3] && FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid);
  end

  assign _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_spinal_port1;
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[0];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_pageFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[1];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_accessFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[2];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[20 : 3];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[40 : 21];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowRead = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[41];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowWrite = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[42];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowExecute = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[43];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowUser = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[44];
  assign _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_spinal_port1;
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[0];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_pageFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[1];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_accessFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[2];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[20 : 3];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[40 : 21];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowRead = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[41];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowWrite = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[42];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowExecute = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[43];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowUser = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[44];
  assign _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_spinal_port1;
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[0];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_pageFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[1];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_accessFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[2];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[20 : 3];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[40 : 21];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowRead = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[41];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowWrite = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[42];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowExecute = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[43];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowUser = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[44];
  assign FetchCachePlugin_logic_translationPort_logic_read_1_readAddress = FetchPlugin_stages_1_Fetch_FETCH_PC[23 : 22];
  assign _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid = FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_spinal_port1;
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[0];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_pageFault = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[1];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_accessFault = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[2];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[10 : 3];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[20 : 11];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowRead = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[21];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowWrite = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[22];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowExecute = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[23];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowUser = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[24];
  always @(*) begin
    FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID[0] = (FetchPlugin_stages_1_MMU_L1_ENTRIES_0_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 24]);
    FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID[1] = (FetchPlugin_stages_1_MMU_L1_ENTRIES_1_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 24]);
  end

  always @(*) begin
    FetchPlugin_stages_1_MMU_L1_HITS[0] = (FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID[0] && FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid);
    FetchPlugin_stages_1_MMU_L1_HITS[1] = (FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID[1] && FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid);
  end

  assign _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid = FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_spinal_port1;
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[0];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_pageFault = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[1];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_accessFault = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[2];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[10 : 3];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[20 : 11];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowRead = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[21];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowWrite = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[22];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowExecute = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[23];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowUser = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[24];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits = {FetchPlugin_stages_1_MMU_L1_HITS,FetchPlugin_stages_1_MMU_L0_HITS};
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hit = (|FetchCachePlugin_logic_translationPort_logic_ctrl_hits);
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0 = FetchCachePlugin_logic_translationPort_logic_ctrl_hits;
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[1];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[2];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[3];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_4 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[4];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_5 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[5];
  always @(*) begin
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[0] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[1] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[2] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_1));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[3] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_2));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[4] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_4 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_3));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[5] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_5 && (! (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_4 || FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_3)));
  end

  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_1 = (|{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0});
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_2 = (|{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0}});
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_3 = (|{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0}}});
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_oh = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[1];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[2];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[3];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[4];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[5];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_6[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineException = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineException[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated : _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_2) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_3 : _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_5)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_6 : _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_8) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_9 : _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_11))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_12 : 32'h00000000) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_13 : 32'h00000000)));
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault[0];
  always @(*) begin
    FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup = (MmuPlugin_logic_satp_mode == 1'b1);
    if(when_MmuPlugin_l315_1) begin
      FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
    if(when_MmuPlugin_l316_1) begin
      FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
  end

  assign FetchCachePlugin_logic_translationPort_logic_ctrl_needRefill = ((FetchPlugin_stages_1_valid && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hit)) && FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup);
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_askRefill = (FetchCachePlugin_logic_translationPort_logic_ctrl_needRefill && FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded);
  assign when_MmuPlugin_l315_1 = ((! MmuPlugin_logic_status_mprv) && (PrivilegedPlugin_setup_privilege == 2'b11));
  assign when_MmuPlugin_l316_1 = (PrivilegedPlugin_setup_privilege == 2'b11);
  assign FetchPlugin_stages_1_MMU_IO = ((ioStartAddr <= FetchPlugin_stages_1_MMU_TRANSLATED) && (FetchPlugin_stages_1_MMU_TRANSLATED <= _zz_FetchPlugin_stages_1_MMU_IO));
  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_REDO = (! FetchCachePlugin_logic_translationPort_logic_ctrl_hit);
    end else begin
      FetchPlugin_stages_1_MMU_REDO = 1'b0;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_TRANSLATED = FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated;
    end else begin
      FetchPlugin_stages_1_MMU_TRANSLATED = FetchPlugin_stages_1_Fetch_FETCH_PC;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_ALLOW_EXECUTE = (FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute && (! (FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser && (PrivilegedPlugin_setup_privilege == 2'b01))));
    end else begin
      FetchPlugin_stages_1_MMU_ALLOW_EXECUTE = 1'b1;
    end
    if(when_MmuPlugin_l356_1) begin
      FetchPlugin_stages_1_MMU_ALLOW_EXECUTE = 1'b0;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_ALLOW_READ = (FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      FetchPlugin_stages_1_MMU_ALLOW_READ = 1'b1;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_ALLOW_WRITE = FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      FetchPlugin_stages_1_MMU_ALLOW_WRITE = 1'b1;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_PAGE_FAULT = ((FetchCachePlugin_logic_translationPort_logic_ctrl_lineException || ((FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser && (PrivilegedPlugin_setup_privilege == 2'b01)) && (! MmuPlugin_logic_status_sum))) || ((! FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser) && (PrivilegedPlugin_setup_privilege == 2'b00)));
    end else begin
      FetchPlugin_stages_1_MMU_PAGE_FAULT = 1'b0;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_ACCESS_FAULT = FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault;
    end else begin
      FetchPlugin_stages_1_MMU_ACCESS_FAULT = (1'b0 || (! (1'b1 || FetchPlugin_stages_1_MMU_IO)));
    end
  end

  assign when_MmuPlugin_l356_1 = (! 1'b1);
  assign FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION = (! FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup);
  assign FetchPlugin_stages_1_MMU_WAYS_OH = FetchCachePlugin_logic_translationPort_logic_ctrl_oh;
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_0_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_1_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_2_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_3_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4 = {FetchPlugin_stages_1_MMU_L1_ENTRIES_0_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[21 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5 = {FetchPlugin_stages_1_MMU_L1_ENTRIES_1_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[21 : 0]};
  assign MmuPlugin_logic_refill_wantExit = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_wantStart = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
        MmuPlugin_logic_refill_wantStart = 1'b1;
      end
    endcase
  end

  assign MmuPlugin_logic_refill_wantKill = 1'b0;
  assign MmuPlugin_logic_refill_busy = (! (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_enumDef_IDLE));
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask = MmuPlugin_logic_refill_portOhReg[0];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask = MmuPlugin_logic_refill_portOhReg[1];
  assign MmuPlugin_logic_refill_portsRequests = {FetchCachePlugin_logic_translationPort_logic_ctrl_askRefill,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_askRefill};
  always @(*) begin
    MmuPlugin_logic_refill_portsRequest = (|MmuPlugin_logic_refill_portsRequests);
    if(when_MmuPlugin_l522) begin
      MmuPlugin_logic_refill_portsRequest = 1'b0;
    end
    if(when_MmuPlugin_l535) begin
      MmuPlugin_logic_refill_portsRequest = 1'b0;
    end
  end

  assign MmuPlugin_logic_refill_portsRequests_ohFirst_input = MmuPlugin_logic_refill_portsRequests;
  assign MmuPlugin_logic_refill_portsRequests_ohFirst_masked = (MmuPlugin_logic_refill_portsRequests_ohFirst_input & (~ _zz_MmuPlugin_logic_refill_portsRequests_ohFirst_masked));
  assign MmuPlugin_logic_refill_portsOh = MmuPlugin_logic_refill_portsRequests_ohFirst_masked;
  assign MmuPlugin_logic_refill_portsAddress = ((MmuPlugin_logic_refill_portsOh_regNext[0] ? _zz_MmuPlugin_logic_refill_portsAddress : 32'h00000000) | (MmuPlugin_logic_refill_portsOh_regNext[1] ? _zz_MmuPlugin_logic_refill_portsAddress_1 : 32'h00000000));
  always @(*) begin
    MmuPlugin_logic_refill_cacheRefillSet = 2'b00;
    if(when_MmuPlugin_l418) begin
      MmuPlugin_logic_refill_cacheRefillSet = MmuPlugin_setup_cacheLoad_rsp_payload_refillSlot;
    end
  end

  always @(*) begin
    MmuPlugin_logic_refill_cacheRefillAnySet = 1'b0;
    if(when_MmuPlugin_l418) begin
      MmuPlugin_logic_refill_cacheRefillAnySet = MmuPlugin_setup_cacheLoad_rsp_payload_refillSlotAny;
    end
  end

  assign FetchCachePlugin_logic_translationPort_wake = MmuPlugin_logic_refill_doWake;
  assign Lsu2Plugin_logic_sharedPip_translationPort_wake = MmuPlugin_logic_refill_doWake;
  assign MmuPlugin_logic_refill_load_readed = MmuPlugin_logic_refill_load_rsp_payload_data[31 : 0];
  assign when_MmuPlugin_l418 = (MmuPlugin_setup_cacheLoad_rsp_valid && MmuPlugin_setup_cacheLoad_rsp_payload_redo);
  always @(*) begin
    MmuPlugin_setup_cacheLoad_cmd_valid = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
        if(when_MmuPlugin_l482) begin
          MmuPlugin_setup_cacheLoad_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
        if(when_MmuPlugin_l482_1) begin
          MmuPlugin_setup_cacheLoad_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_setup_cacheLoad_cmd_payload_virtual = MmuPlugin_logic_refill_load_address;
  assign MmuPlugin_setup_cacheLoad_cmd_payload_size = 2'b10;
  assign MmuPlugin_setup_cacheLoad_cmd_payload_redoOnDataHazard = 1'b1;
  assign MmuPlugin_setup_cacheLoad_cmd_payload_unlocked = 1'b0;
  assign MmuPlugin_setup_cacheLoad_cmd_payload_unique = 1'b0;
  assign MmuPlugin_setup_cacheLoad_translated_physical = MmuPlugin_logic_refill_load_address;
  assign MmuPlugin_setup_cacheLoad_translated_abord = 1'b0;
  assign MmuPlugin_setup_cacheLoad_cancels = 3'b000;
  assign _zz_MmuPlugin_logic_refill_load_flags_V = MmuPlugin_logic_refill_load_readed;
  assign MmuPlugin_logic_refill_load_flags_V = _zz_MmuPlugin_logic_refill_load_flags_V[0];
  assign MmuPlugin_logic_refill_load_flags_R = _zz_MmuPlugin_logic_refill_load_flags_V[1];
  assign MmuPlugin_logic_refill_load_flags_W = _zz_MmuPlugin_logic_refill_load_flags_V[2];
  assign MmuPlugin_logic_refill_load_flags_X = _zz_MmuPlugin_logic_refill_load_flags_V[3];
  assign MmuPlugin_logic_refill_load_flags_U = _zz_MmuPlugin_logic_refill_load_flags_V[4];
  assign MmuPlugin_logic_refill_load_flags_G = _zz_MmuPlugin_logic_refill_load_flags_V[5];
  assign MmuPlugin_logic_refill_load_flags_A = _zz_MmuPlugin_logic_refill_load_flags_V[6];
  assign MmuPlugin_logic_refill_load_flags_D = _zz_MmuPlugin_logic_refill_load_flags_V[7];
  assign MmuPlugin_logic_refill_load_leaf = (MmuPlugin_logic_refill_load_flags_R || MmuPlugin_logic_refill_load_flags_X);
  always @(*) begin
    MmuPlugin_logic_refill_load_exception = ((((! MmuPlugin_logic_refill_load_flags_V) || ((! MmuPlugin_logic_refill_load_flags_R) && MmuPlugin_logic_refill_load_flags_W)) || MmuPlugin_logic_refill_load_rsp_payload_fault) || ((! MmuPlugin_logic_refill_load_leaf) && ((MmuPlugin_logic_refill_load_flags_D || MmuPlugin_logic_refill_load_flags_A) || MmuPlugin_logic_refill_load_flags_U)));
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(when_MmuPlugin_l491) begin
          MmuPlugin_logic_refill_load_exception = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_load_levelException_0 = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_load_levelException_1 = 1'b0;
    if(when_MmuPlugin_l446) begin
      MmuPlugin_logic_refill_load_levelException_1 = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_nextLevelBase = 32'h00000000;
    MmuPlugin_logic_refill_load_nextLevelBase[21 : 12] = MmuPlugin_logic_refill_load_readed[19 : 10];
    MmuPlugin_logic_refill_load_nextLevelBase[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 = 32'h00000000;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[21 : 12] = MmuPlugin_logic_refill_load_readed[19 : 10];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 = 32'h00000000;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[21 : 12] = MmuPlugin_logic_refill_virtual[21 : 12];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  assign when_MmuPlugin_l446 = (MmuPlugin_logic_refill_load_readed[19 : 10] != 10'h000);
  always @(*) begin
    MmuPlugin_logic_invalidate_canStart = 1'b1;
    if(when_MmuPlugin_l541) begin
      MmuPlugin_logic_invalidate_canStart = 1'b0;
    end
  end

  assign MmuPlugin_logic_invalidate_done = MmuPlugin_logic_invalidate_counter[2];
  assign when_MmuPlugin_l522 = (! MmuPlugin_logic_invalidate_done);
  assign FetchPlugin_stages_0_haltRequest_MmuPlugin_l533 = ((! MmuPlugin_logic_invalidate_done) || MmuPlugin_logic_invalidate_requested);
  assign when_MmuPlugin_l535 = (MmuPlugin_logic_invalidate_requested && MmuPlugin_logic_invalidate_canStart);
  assign when_MmuPlugin_l541 = (MmuPlugin_logic_refill_busy || (|Lsu2Plugin_setup_postCommitBusy));
  assign when_MmuPlugin_l545 = (MmuPlugin_logic_invalidate_done && (! MmuPlugin_logic_invalidate_done_regNext));
  assign Lsu2Plugin_logic_sharedPip_stages_3_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_2_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_1_isRemoved = (Lsu2Plugin_logic_sharedPip_stages_1_isFlushed || Lsu2Plugin_logic_sharedPip_stages_1_isThrown);
  assign Lsu2Plugin_logic_sharedPip_stages_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_1_isThrown = 1'b0;
  assign Lsu2Plugin_logic_sharedPip_stages_0_isRemoved = (Lsu2Plugin_logic_sharedPip_stages_0_isFlushed || Lsu2Plugin_logic_sharedPip_stages_0_isThrown);
  assign Lsu2Plugin_logic_sharedPip_stages_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_0_isThrown = 1'b0;
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_valid = Lsu2Plugin_logic_sharedPip_stages_0_valid;
    if(when_Pipeline_l278) begin
      _zz_Lsu2Plugin_logic_sharedPip_stages_1_valid = 1'b0;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_ready = 1'b1;
    if(when_Pipeline_l278) begin
      Lsu2Plugin_logic_sharedPip_stages_0_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278 = (|Lsu2Plugin_logic_sharedPip_stages_0_haltRequest_Lsu2Plugin_l990);
  assign Lsu2Plugin_logic_sharedPip_stages_1_ready = 1'b1;
  assign Lsu2Plugin_logic_sharedPip_stages_2_ready = 1'b1;
  assign Lsu2Plugin_logic_sharedPip_stages_3_ready = 1'b1;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_valid = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_data = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_data;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_fault = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_fault;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_redo = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_redo;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlot = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlot;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlotAny = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_resulting = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
  assign Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_resulting = Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_overloaded;
  assign Lsu2Plugin_logic_lqSqArbitration_s1_isRemoved = (Lsu2Plugin_logic_lqSqArbitration_s1_isFlushed || Lsu2Plugin_logic_lqSqArbitration_s1_isThrown);
  assign Lsu2Plugin_logic_lqSqArbitration_s1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_lqSqArbitration_s1_isThrown = 1'b0;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_ready = Lsu2Plugin_logic_lqSqArbitration_s0_ready_output;
  always @(*) begin
    Lsu2Plugin_logic_lqSqArbitration_s1_ready = 1'b1;
    if(when_Pipeline_l278_1) begin
      Lsu2Plugin_logic_lqSqArbitration_s1_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_1 = (|{Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842,Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l834});
  always @(*) begin
    Lsu2Plugin_logic_lqSqArbitration_s0_ready_output = Lsu2Plugin_logic_lqSqArbitration_s1_ready;
    if(when_Connection_l74) begin
      Lsu2Plugin_logic_lqSqArbitration_s0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74 = (! Lsu2Plugin_logic_lqSqArbitration_s1_valid);
  always @(*) begin
    Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_stateReg;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
        if(when_Lsu2Plugin_l1704) begin
          if(when_Lsu2Plugin_l1705) begin
            Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY;
          end
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
        if(Lsu2Plugin_setup_cacheLoad_cmd_fire) begin
          Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP;
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
        if(Lsu2Plugin_setup_cacheLoad_rsp_valid) begin
          if(Lsu2Plugin_setup_cacheLoad_rsp_payload_redo) begin
            Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD;
          end else begin
            if(Lsu2Plugin_setup_cacheLoad_rsp_payload_fault) begin
              Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_TRAP;
            end else begin
              Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_ALU;
            end
          end
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
        if(when_Lsu2Plugin_l1715) begin
          if(Lsu2Plugin_logic_special_storeSc) begin
            Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_ALU;
          end else begin
            Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD;
          end
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
        Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
        Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_SYNC;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
        if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
          Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_IDLE;
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
        Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
        Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_IDLE;
      end
      default : begin
      end
    endcase
    if(Lsu2Plugin_logic_special_atomic_wantStart) begin
      Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_IDLE;
    end
    if(Lsu2Plugin_logic_special_atomic_wantKill) begin
      Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_BOOT;
    end
  end

  assign when_Lsu2Plugin_l1704 = (Lsu2Plugin_logic_special_enabled && Lsu2Plugin_logic_special_isAtomic);
  assign when_Lsu2Plugin_l1705 = (Lsu2Plugin_logic_sq_ptr_commit == Lsu2Plugin_logic_sq_ptr_free);
  assign Lsu2Plugin_setup_cacheLoad_cmd_fire = (Lsu2Plugin_setup_cacheLoad_cmd_valid && Lsu2Plugin_setup_cacheLoad_cmd_ready);
  assign when_Lsu2Plugin_l1715 = (&Lsu2Plugin_logic_special_atomic_lockDelayCounter);
  assign when_Lsu2Plugin_l1828 = (Lsu2Plugin_logic_special_storeSc && (! Lsu2Plugin_logic_special_atomic_gotReservation));
  assign when_StateMachine_l253 = ((! (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID])) && (Lsu2Plugin_logic_special_atomic_stateNext[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]));
  assign when_StateMachine_l253_1 = ((! (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID])) && (Lsu2Plugin_logic_special_atomic_stateNext[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]));
  always @(*) begin
    MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_stateReg;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
        if(MmuPlugin_logic_refill_portsRequest) begin
          MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_INIT;
        end
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
        MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_1;
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
        if(when_MmuPlugin_l482) begin
          if(MmuPlugin_setup_cacheLoad_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_RSP_0;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
        if(when_MmuPlugin_l482_1) begin
          if(MmuPlugin_setup_cacheLoad_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_RSP_1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_0;
          end else begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_1;
          end else begin
            if(when_MmuPlugin_l499) begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
            end else begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_0;
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(MmuPlugin_logic_refill_wantStart) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
    end
    if(MmuPlugin_logic_refill_wantKill) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_BOOT;
    end
  end

  assign when_MmuPlugin_l482 = ((MmuPlugin_logic_refill_cacheRefill == 2'b00) && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l482_1 = ((MmuPlugin_logic_refill_cacheRefill == 2'b00) && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l491 = (! MmuPlugin_logic_refill_load_leaf);
  assign when_MmuPlugin_l499 = (MmuPlugin_logic_refill_load_leaf || MmuPlugin_logic_refill_load_exception);
  assign MmuPlugin_logic_refill_doWake = (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_enumDef_IDLE);
  assign DecoderPlugin_logic_slots_0_rdZero = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[11 : 7] == 5'h00);
  assign FrontendPlugin_decoded_LEGAL_0 = ((|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000005f) == 32'h00000017),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000007f) == 32'h0000006f),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_LEGAL_0) == 32'h00001073),{(_zz_FrontendPlugin_decoded_LEGAL_0_1 == _zz_FrontendPlugin_decoded_LEGAL_0_2),{_zz_FrontendPlugin_decoded_LEGAL_0_3,{_zz_FrontendPlugin_decoded_LEGAL_0_4,_zz_FrontendPlugin_decoded_LEGAL_0_5}}}}}}) && (! FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_0));
  assign FrontendPlugin_decoded_READ_RS_0_0 = _zz_FrontendPlugin_decoded_READ_RS_0_0[0];
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_0 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h10000070) == 32'h00000020);
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_0_1 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h08000070) == 32'h08000020);
  assign FrontendPlugin_decoded_READ_RS_1_0 = _zz_FrontendPlugin_decoded_READ_RS_1_0[0];
  assign _zz_260 = zz_DecoderPlugin_logic_slots_0_x0AlwaysZero(1'b0);
  always @(*) DecoderPlugin_logic_slots_0_x0AlwaysZero = _zz_260;
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000048) == 32'h00000048);
  assign FrontendPlugin_decoded_WRITE_RD_0 = (_zz_FrontendPlugin_decoded_WRITE_RD_0_1[0] && (! (DecoderPlugin_logic_slots_0_rdZero && DecoderPlugin_logic_slots_0_x0AlwaysZero)));
  assign FrontendPlugin_decoded_ALU0_SEL_0 = _zz_FrontendPlugin_decoded_ALU0_SEL_0[0];
  assign FrontendPlugin_decoded_EU0_SEL_0 = _zz_FrontendPlugin_decoded_EU0_SEL_0[0];
  assign FrontendPlugin_decoded_LQ_ALLOC_0 = _zz_FrontendPlugin_decoded_LQ_ALLOC_0[0];
  assign FrontendPlugin_decoded_SQ_ALLOC_0 = _zz_FrontendPlugin_decoded_SQ_ALLOC_0_2[0];
  assign FrontendPlugin_decoded_TRAP_0 = (FrontendPlugin_decoded_Frontend_MASK_ALIGNED_0 && ((((! FrontendPlugin_decoded_LEGAL_0) || FrontendPlugin_decoded_Frontend_FETCH_FAULT_0) || DecoderPlugin_setup_trapRaise) || DecoderPlugin_setup_debugEnter_0));
  assign FrontendPlugin_decoded_Frontend_DECODED_MASK_0 = (FrontendPlugin_decoded_Frontend_MASK_ALIGNED_0 && (! (|FrontendPlugin_decoded_TRAP_0)));
  assign FrontendPlugin_decoded_Frontend_MICRO_OP_0 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0;
  assign FrontendPlugin_decoded_ARCH_RD_0 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[11 : 7];
  assign FrontendPlugin_decoded_ARCH_RS_0_0 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[19 : 15];
  assign FrontendPlugin_decoded_ARCH_RS_1_0 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[24 : 20];
  assign DecoderPlugin_logic_exception_set = (FrontendPlugin_decoded_isFireing && (|FrontendPlugin_decoded_TRAP_0));
  assign DecoderPlugin_logic_exception_clear = FrontendPlugin_decoded_isFlushed;
  assign when_DecoderPlugin_l302 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l303 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l304 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l306 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l307 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l308 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l309 = (! DecoderPlugin_logic_exception_trigged);
  assign DecoderPlugin_logic_exception_compressedFault = _zz_DecoderPlugin_logic_exception_compressedFault[0];
  assign DecoderPlugin_logic_exception_fetchFault = _zz_DecoderPlugin_logic_exception_fetchFault[0];
  assign DecoderPlugin_logic_exception_fetchFaultPage = _zz_DecoderPlugin_logic_exception_fetchFaultPage[0];
  assign DecoderPlugin_logic_exception_debugEnter = _zz_DecoderPlugin_logic_exception_debugEnter[0];
  assign DecoderPlugin_logic_exception_pc = (DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_epcReg_0 : 32'h00000000);
  assign DecoderPlugin_logic_exception_pipelineEmpty = ((! FrontendPlugin_isBusyAfterDecode) && CommitPlugin_setup_isRobEmpty);
  assign DecoderPlugin_logic_exception_doIt = (DecoderPlugin_logic_exception_trigged && DecoderPlugin_logic_exception_pipelineEmpty);
  assign _zz_FrontendPlugin_decoded_isFlushingRoot = (DecoderPlugin_logic_exception_doIt || DecoderPlugin_logic_exception_doItAgain);
  assign FrontendPlugin_decoded_haltRequest_DecoderPlugin_l324 = DecoderPlugin_logic_exception_trigged;
  assign FrontendPlugin_decoded_haltRequest_DecoderPlugin_l325 = (DecoderPlugin_setup_trapHalt && (! DecoderPlugin_setup_trapRaise));
  assign DecoderPlugin_setup_trapReady = (FrontendPlugin_decoded_valid && DecoderPlugin_logic_exception_pipelineEmpty);
  assign DecoderPlugin_setup_exceptionPort_valid = DecoderPlugin_logic_exception_doIt;
  assign DecoderPlugin_setup_exceptionPort_payload_epc = DecoderPlugin_logic_exception_pc;
  always @(*) begin
    if(DecoderPlugin_logic_exception_fetchFault) begin
      if(DecoderPlugin_logic_exception_fetchFaultPage) begin
        DecoderPlugin_setup_exceptionPort_payload_cause = 4'b1100;
      end else begin
        DecoderPlugin_setup_exceptionPort_payload_cause = 4'b0001;
      end
    end else begin
      if(DecoderPlugin_logic_exception_compressedFault) begin
        DecoderPlugin_setup_exceptionPort_payload_cause = 4'b0010;
      end else begin
        DecoderPlugin_setup_exceptionPort_payload_cause = 4'b0010;
      end
    end
  end

  always @(*) begin
    if(DecoderPlugin_logic_exception_fetchFault) begin
      DecoderPlugin_setup_exceptionPort_payload_tval = _zz_DecoderPlugin_setup_exceptionPort_payload_tval;
    end else begin
      if(DecoderPlugin_logic_exception_compressedFault) begin
        DecoderPlugin_setup_exceptionPort_payload_tval = ((DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_instReg_0 : 32'h00000000) & 32'h0000ffff);
      end else begin
        DecoderPlugin_setup_exceptionPort_payload_tval = (DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_instReg_0 : 32'h00000000);
      end
    end
  end

  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h00001048) == 32'h00001008);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_1 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h00002050) == 32'h00002050);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_2 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h02000050) == 32'h02000050);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_3 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h00001050) == 32'h00001050);
  assign FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0[0];
  assign FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0[0];
  assign FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_4[0];
  assign FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0[0];
  assign FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0[0];
  assign FrontendPlugin_dispatch_LATENCY_0_0 = (|{((FrontendPlugin_dispatch_Frontend_MICRO_OP_0 & 32'h00000030) == 32'h00000010),{((FrontendPlugin_dispatch_Frontend_MICRO_OP_0 & 32'h0000004c) == 32'h00000004),((FrontendPlugin_dispatch_Frontend_MICRO_OP_0 & 32'h02000050) == 32'h00000010)}});
  assign FrontendPlugin_decoded_IS_JAL_0 = _zz_FrontendPlugin_decoded_IS_JAL_0[0];
  assign FrontendPlugin_decoded_IS_JALR_0 = _zz_FrontendPlugin_decoded_IS_JALR_0[0];
  assign FrontendPlugin_decoded_Prediction_IS_BRANCH_0 = _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_0[0];
  assign FrontendPlugin_decoded_IS_ANY_0 = _zz_FrontendPlugin_decoded_IS_ANY_0[0];
  assign switch_Misc_l241_2 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[2];
  always @(*) begin
    case(switch_Misc_l241_2)
      1'b0 : begin
        _zz_FrontendPlugin_decoded_OFFSET_0 = {{19{_zz__zz_FrontendPlugin_decoded_OFFSET_0[12]}}, _zz__zz_FrontendPlugin_decoded_OFFSET_0};
      end
      default : begin
        _zz_FrontendPlugin_decoded_OFFSET_0 = {{11{_zz__zz_FrontendPlugin_decoded_OFFSET_0_1[20]}}, _zz__zz_FrontendPlugin_decoded_OFFSET_0_1};
      end
    endcase
  end

  assign FrontendPlugin_decoded_OFFSET_0 = _zz_FrontendPlugin_decoded_OFFSET_0;
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink = (|{(FrontendPlugin_decoded_ARCH_RD_0 == 5'h05),(FrontendPlugin_decoded_ARCH_RD_0 == 5'h01)});
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rs1Link = (|{(FrontendPlugin_decoded_ARCH_RS_0_0 == 5'h05),(FrontendPlugin_decoded_ARCH_RS_0_0 == 5'h01)});
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdEquRs1 = (FrontendPlugin_decoded_ARCH_RD_0 == FrontendPlugin_decoded_ARCH_RS_0_0);
  assign FrontendPlugin_decoded_RAS_PUSH_0 = ((FrontendPlugin_decoded_IS_JAL_0 || FrontendPlugin_decoded_IS_JALR_0) && DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink);
  assign FrontendPlugin_decoded_RAS_POP_0 = (FrontendPlugin_decoded_IS_JALR_0 && (((! DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink) && DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rs1Link) || ((DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink && DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rs1Link) && (! DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdEquRs1))));
  assign FrontendPlugin_decoded_CONDITIONAL_PREDICTION_0 = FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_0[0];
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices = (_zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices + {1'b0,1'b1});
  assign FrontendPlugin_decoded_PC_INC_0 = _zz_FrontendPlugin_decoded_PC_INC_0;
  assign FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0 = ($signed(_zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0) + $signed(FrontendPlugin_decoded_OFFSET_0));
  assign FrontendPlugin_decoded_BAD_RET_PC_0 = (FrontendPlugin_decoded_RAS_POP_0 && (DecoderPredictionPlugin_logic_ras_read != FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_0));
  assign FrontendPlugin_decoded_CAN_IMPROVE_0 = ((! FrontendPlugin_decoded_IS_JALR_0) || FrontendPlugin_decoded_RAS_POP_0);
  assign FrontendPlugin_decoded_BRANCHED_PREDICTION_0 = (((FrontendPlugin_decoded_Prediction_IS_BRANCH_0 && FrontendPlugin_decoded_CONDITIONAL_PREDICTION_0) || FrontendPlugin_decoded_IS_JAL_0) || FrontendPlugin_decoded_IS_JALR_0);
  always @(*) begin
    FrontendPlugin_serialized_PC_TARGET_0 = FrontendPlugin_serialized_PC_TARGET_PRE_RAS_0;
    if(FrontendPlugin_serialized_IS_JALR_0) begin
      FrontendPlugin_serialized_PC_TARGET_0 = DecoderPredictionPlugin_logic_ras_read;
    end
  end

  assign FrontendPlugin_serialized_PC_PREDICTION_0 = (FrontendPlugin_serialized_BRANCHED_PREDICTION_0 ? FrontendPlugin_serialized_PC_TARGET_0 : FrontendPlugin_serialized_PC_INC_0);
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_applyIt_badTaken = (FrontendPlugin_serialized_IS_ANY_0 ? (FrontendPlugin_serialized_BRANCHED_PREDICTION_0 != FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0) : FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0);
  assign FrontendPlugin_serialized_MISSMATCH_PC_0 = (DecoderPredictionPlugin_logic_decodePatch_slots_0_applyIt_badTaken || FrontendPlugin_serialized_BAD_RET_PC_0);
  assign FrontendPlugin_serialized_MISSMATCH_HISTORY_0 = 1'b0;
  assign FrontendPlugin_serialized_MISSMATCH_0 = (FrontendPlugin_serialized_MISSMATCH_PC_0 || FrontendPlugin_serialized_MISSMATCH_HISTORY_0);
  assign FrontendPlugin_serialized_NEED_CORRECTION_0 = ((FrontendPlugin_serialized_Frontend_DECODED_MASK_0 && FrontendPlugin_serialized_CAN_IMPROVE_0) && FrontendPlugin_serialized_MISSMATCH_0);
  assign FrontendPlugin_serialized_BRANCH_SEL_0 = FrontendPlugin_serialized_IS_ANY_0;
  always @(*) begin
    if(FrontendPlugin_serialized_NEED_CORRECTION_0) begin
      FrontendPlugin_serialized_BRANCH_EARLY_0_taken = FrontendPlugin_serialized_BRANCHED_PREDICTION_0;
    end else begin
      FrontendPlugin_serialized_BRANCH_EARLY_0_taken = FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0;
    end
  end

  always @(*) begin
    if(FrontendPlugin_serialized_NEED_CORRECTION_0) begin
      FrontendPlugin_serialized_BRANCH_EARLY_0_pc = FrontendPlugin_serialized_PC_TARGET_0;
    end else begin
      FrontendPlugin_serialized_BRANCH_EARLY_0_pc = FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
    end
  end

  assign when_DecoderPredictionPlugin_l212 = (FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0 && FrontendPlugin_serialized_RAS_PUSH_0);
  assign when_DecoderPredictionPlugin_l213 = (! DecoderPredictionPlugin_logic_decodePatch_rasPushUsed);
  assign when_DecoderPredictionPlugin_l219 = (FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0 && FrontendPlugin_serialized_RAS_POP_0);
  assign FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_0 = DecoderPredictionPlugin_logic_ras_ptr_push;
  assign DecoderPredictionPlugin_logic_decodePatch_applyIt_hit = (|FrontendPlugin_serialized_NEED_CORRECTION_0);
  assign FrontendPlugin_serialized_isFireing = (FrontendPlugin_serialized_valid && FrontendPlugin_serialized_ready);
  assign when_DecoderPredictionPlugin_l236 = (FrontendPlugin_serialized_ready || FrontendPlugin_serialized_isFlushed);
  assign DecoderPredictionPlugin_setup_decodeJump_valid = (FrontendPlugin_serialized_valid && DecoderPredictionPlugin_logic_decodePatch_applyIt_hit);
  assign DecoderPredictionPlugin_setup_decodeJump_payload_pc = FrontendPlugin_serialized_PC_PREDICTION_0;
  assign DecoderPredictionPlugin_setup_historyPush_flush = DecoderPredictionPlugin_setup_decodeJump_valid;
  assign when_DecoderPredictionPlugin_l243 = (! FrontendPlugin_serialized_isFireing);
  assign when_DecoderPredictionPlugin_l244 = (! FrontendPlugin_serialized_isFireing);
  assign FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0 = (FrontendPlugin_serialized_Frontend_DECODED_MASK_0 && (! 1'b0));
  assign DecoderPredictionPlugin_setup_historyPush_mask[0] = ((((FrontendPlugin_serialized_valid && DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle) && FrontendPlugin_serialized_Prediction_IS_BRANCH_0) && FrontendPlugin_serialized_Frontend_DECODED_MASK_0) && (! 1'b0));
  assign DecoderPredictionPlugin_setup_historyPush_taken[0] = FrontendPlugin_serialized_BRANCHED_PREDICTION_0;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_valid = ALU0_ExecutionUnitBase_pipeline_push_port_valid;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID = ALU0_ExecutionUnitBase_pipeline_push_port_robId;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD = ALU0_ExecutionUnitBase_pipeline_push_port_physRd;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1[31 : 0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1[5 : 0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1[5 : 0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_PC = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_1[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL = ((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000004) == 32'h00000004);
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1 = {(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004004) == 32'h00004000)),(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00006004) == 32'h00002000))};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED = ((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001000) == 32'h00001000);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1 = {(|_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED),(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00003000) == 32'h00002000))};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL = (|_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL);
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL = {(|_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL),(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000024) == 32'h00000000))};
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid = ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  assign ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address = ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1 = ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  assign ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid = ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  assign ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address = ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2 = ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  assign ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid = ((ALU0_ExecutionUnitBase_pipeline_execute_0_valid && ALU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD) && (|ALU0_IntFormatPlugin_logic_stages_0_wb_valid));
  assign ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId = ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_address = ALU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  assign ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_data = ALU0_IntFormatPlugin_logic_stages_0_wb_payload;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_isFireing = (ALU0_ExecutionUnitBase_pipeline_execute_0_valid && ALU0_ExecutionUnitBase_pipeline_execute_0_ready);
  assign ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid = (ALU0_ExecutionUnitBase_pipeline_execute_0_isFireing && ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0);
  assign ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id = ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ready = 1'b1;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_valid = ALU0_ExecutionUnitBase_pipeline_fetch_1_valid;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2 = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL = ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL = ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL = ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL = ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT = ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED = ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD = ALU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID = ALU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD = ALU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0 = ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_valid = EU0_ExecutionUnitBase_pipeline_push_port_valid;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID = EU0_ExecutionUnitBase_pipeline_push_port_robId;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD = EU0_ExecutionUnitBase_pipeline_push_port_physRd;
  assign EU0_ExecutionUnitBase_pipeline_push_port_ready = EU0_ExecutionUnitBase_pipeline_fetch_0_ready;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0 = EU0_ExecutionUnitBase_pipeline_push_port_context_0;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1 = EU0_ExecutionUnitBase_pipeline_push_port_context_1;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1[31 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_PC = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_1[31 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1[1 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_1[3 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_1[0 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000040) == 32'h00000040);
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002000) == 32'h00002000);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001000) == 32'h00001000);
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00006000) == 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000008) == 32'h00000008);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1 = {(|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h0000000c) == 32'h00000004)),(|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO)};
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000020) == 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL = {(|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD),(|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000060) == 32'h00000020))};
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1[0];
  assign EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid = EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  assign EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address = EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1 = EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  assign EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid = EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  assign EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address = EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2 = EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid = ((EU0_ExecutionUnitBase_pipeline_execute_2_valid && EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD) && (|EU0_IntFormatPlugin_logic_stages_0_wb_valid));
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_address = EU0_ExecutionUnitBase_pipeline_execute_2_PHYS_RD;
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_data = EU0_IntFormatPlugin_logic_stages_0_wb_payload;
  assign EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_ExecutionUnitBase_l303 = (EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid && (! EU0_ExecutionUnitBase_pipeline_writeBack_0_write_ready));
  assign EU0_ExecutionUnitBase_pipeline_completion_0_port_valid = (EU0_ExecutionUnitBase_pipeline_execute_2_isFireing && EU0_ExecutionUnitBase_pipeline_execute_2_completion_SEL_E2);
  assign EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_fire = (EU0_ExecutionUnitBase_pipeline_execute_2_isFireing && (|{EU0_CsrAccessPlugin_logic_wake_wakeRobsSel,{EU0_BranchPlugin_logic_wake_wakeRobsSel,{EU0_DivPlugin_logic_wake_wakeRobsSel,EU0_MulPlugin_logic_wake_wakeRobsSel}}}));
  assign EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_valid = (EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_fire && EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD);
  assign EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_fire = (EU0_ExecutionUnitBase_pipeline_execute_2_isFireing && (|{EU0_CsrAccessPlugin_logic_wake_wakeRegFileSel,{EU0_BranchPlugin_logic_wake_wakeRegFileSel,{EU0_DivPlugin_logic_wake_wakeRegFileSel,EU0_MulPlugin_logic_wake_wakeRegFileSel}}}));
  assign EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_valid = (EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_fire && EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD);
  assign EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_payload_physical = EU0_ExecutionUnitBase_pipeline_execute_2_PHYS_RD;
  assign EU0_ExecutionUnitBase_pipeline_execute_2_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_execute_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_isRemoved = (EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed || EU0_ExecutionUnitBase_pipeline_execute_0_isThrown);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_isThrown = 1'b0;
  assign EU0_ExecutionUnitBase_pipeline_fetch_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_ready = EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output;
  assign EU0_ExecutionUnitBase_pipeline_fetch_1_ready = EU0_ExecutionUnitBase_pipeline_fetch_1_ready_output;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_valid = EU0_ExecutionUnitBase_pipeline_execute_0_valid;
    if(when_Pipeline_l278_2) begin
      _zz_EU0_ExecutionUnitBase_pipeline_execute_1_valid = 1'b0;
    end
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_0_ready = EU0_ExecutionUnitBase_pipeline_execute_0_ready_output;
    if(when_Pipeline_l278_2) begin
      EU0_ExecutionUnitBase_pipeline_execute_0_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_2 = (|EU0_ExecutionUnitBase_pipeline_execute_0_haltRequest_DivPlugin_l83);
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_valid = EU0_ExecutionUnitBase_pipeline_execute_1_valid;
    if(when_Pipeline_l278_3) begin
      _zz_EU0_ExecutionUnitBase_pipeline_execute_2_valid = 1'b0;
    end
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_1_ready = EU0_ExecutionUnitBase_pipeline_execute_1_ready_output;
    if(when_Pipeline_l278_3) begin
      EU0_ExecutionUnitBase_pipeline_execute_1_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_3 = (|EU0_ExecutionUnitBase_pipeline_execute_1_haltRequest_DivPlugin_l91);
  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_2_ready = 1'b1;
    if(when_Pipeline_l278_4) begin
      EU0_ExecutionUnitBase_pipeline_execute_2_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_4 = (|{EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_ExecutionUnitBase_l303,EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_CsrAccessPlugin_l375});
  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output = EU0_ExecutionUnitBase_pipeline_fetch_1_ready;
    if(when_Connection_l74_1) begin
      EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_1 = (! EU0_ExecutionUnitBase_pipeline_fetch_1_valid);
  assign EU0_ExecutionUnitBase_pipeline_fetch_1_ready_output = EU0_ExecutionUnitBase_pipeline_execute_0_ready;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_valid = EU0_ExecutionUnitBase_pipeline_fetch_1_valid;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2 = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1 = EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS1;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2 = EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS2;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_SIGNED = EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS1_SIGNED;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED = EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS2_SIGNED;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM = EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_REM;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL = EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP = EU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_PC = EU0_ExecutionUnitBase_pipeline_fetch_1_PC;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID = EU0_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID = EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_ROB_MSB = EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_MSB;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SC = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SC;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_AMO = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_AMO;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD = EU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD = EU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_LSU_ID = EU0_ExecutionUnitBase_pipeline_fetch_1_LSU_ID;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LR = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LR;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LOAD = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LOAD;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_IMM = EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_IMM;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK = EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_MASK;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_CLEAR = EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_CLEAR;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_HIGH = EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_HIGH;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_EBREAK = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_EBREAK;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_ECALL = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_ECALL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_XRET = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_XRET;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_I = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_I;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FLUSH_DATA = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FLUSH_DATA;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_VMA = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_VMA;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_WFI = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_WFI;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E2 = EU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E2;
  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_0_ready_output = EU0_ExecutionUnitBase_pipeline_execute_1_ready;
    if(when_Connection_l74_2) begin
      EU0_ExecutionUnitBase_pipeline_execute_0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_2 = (! EU0_ExecutionUnitBase_pipeline_execute_1_valid);
  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_1_ready_output = EU0_ExecutionUnitBase_pipeline_execute_2_ready;
    if(when_Connection_l74_3) begin
      EU0_ExecutionUnitBase_pipeline_execute_1_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_3 = (! EU0_ExecutionUnitBase_pipeline_execute_2_valid);
  assign BranchContextPlugin_free_dispatchMem_writes_0_port_valid = ((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_BRANCH_SEL_0) && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0);
  assign BranchContextPlugin_free_dispatchMem_writes_0_port_payload_address = FrontendPlugin_dispatch_BRANCH_ID_0;
  assign BranchContextPlugin_free_dispatchMem_writes_0_port_payload_data = {FrontendPlugin_dispatch_Prediction_IS_BRANCH_0,{FrontendPlugin_dispatch_GSHARE_COUNTER_0_0,FrontendPlugin_dispatch_BRANCH_HISTORY_0}};
  assign BranchContextPlugin_free_learn_valid = (BranchContextPlugin_logic_ptr_free != BranchContextPlugin_logic_ptr_commited);
  assign BranchContextPlugin_free_learn_bid = BranchContextPlugin_logic_ptr_free[1:0];
  assign _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice = BranchContextPlugin_logic_mem_finalBranch_spinal_port1;
  assign BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice = _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[31 : 0];
  assign BranchContextPlugin_learn_BRANCH_FINAL_pcTarget = _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[63 : 32];
  assign BranchContextPlugin_learn_BRANCH_FINAL_taken = _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[64];
  assign BranchContextPlugin_free_learn_raw = BranchContextPlugin_free_dispatchMem_mem_spinal_port1;
  assign BranchContextPlugin_free_learn_BRANCH_HISTORY = BranchContextPlugin_free_learn_raw[23 : 0];
  assign BranchContextPlugin_free_learn_GSHARE_COUNTER_0 = _zz_BranchContextPlugin_free_learn_GSHARE_COUNTER_0[1 : 0];
  assign BranchContextPlugin_free_learn_Prediction_IS_BRANCH = BranchContextPlugin_free_learn_raw[26];
  assign BranchContextPlugin_setup_learnValid = BranchContextPlugin_free_learn_valid;
  assign DispatchPlugin_logic_queueStaticWakeTransposed_0 = {DispatchPlugin_logic_queue_io_contexts_7_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_6_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_5_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_4_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_3_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_2_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_1_staticWake[0],DispatchPlugin_logic_queue_io_contexts_0_staticWake[0]}}}}}}};
  assign DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0 = DispatchPlugin_logic_queueStaticWakeTransposed_0;
  assign toplevel_DispatchPlugin_logic_queue_io_push_fire = (FrontendPlugin_dispatch_isFireing && DispatchPlugin_logic_queue_io_push_ready);
  assign FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l187 = (! DispatchPlugin_logic_queue_io_push_ready);
  assign DispatchPlugin_logic_push_skip = (! (|FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0));
  assign DispatchPlugin_logic_push_fenceOlder = (FrontendPlugin_dispatch_valid && (|(FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 && FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_0)));
  assign DispatchPlugin_logic_push_fenceYounger = (FrontendPlugin_dispatch_valid && (|(FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 && FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_0)));
  assign when_DispatchPlugin_l192 = (FrontendPlugin_dispatch_isFireing && (! DispatchPlugin_logic_push_skip));
  assign DispatchPlugin_logic_push_commitNotWaitingOnUs = (|(CommitPlugin_logic_commit_head ^ FrontendPlugin_dispatch_ROB_ID));
  assign FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l195 = (DispatchPlugin_logic_push_fenceOlder && DispatchPlugin_logic_push_commitNotWaitingOnUs);
  assign FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l196 = ((DispatchPlugin_logic_push_fenceYoungerLast && DispatchPlugin_logic_push_commitNotWaitingOnUs) && (! DispatchPlugin_logic_push_skip));
  assign DispatchPlugin_logic_push_slots_0_self = ((FrontendPlugin_dispatch_WRITE_RD_0 && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) ? 8'h80 : 8'h00);
  assign DispatchPlugin_logic_push_slots_0_events_0 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_0 ? _zz_DispatchPlugin_logic_push_slots_0_events_0 : 8'h00);
  assign DispatchPlugin_logic_push_slots_0_events_1 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_0 ? _zz_DispatchPlugin_logic_push_slots_0_events_1 : 8'h00);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_0_event = ((DispatchPlugin_logic_push_slots_0_self | DispatchPlugin_logic_push_slots_0_events_0) | DispatchPlugin_logic_push_slots_0_events_1);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_0_sel = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 ? {FrontendPlugin_dispatch_EU0_SEL_0,FrontendPlugin_dispatch_ALU0_SEL_0} : 2'b00);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_0_context_robId = (FrontendPlugin_dispatch_ROB_ID | 4'b0000);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_0_context_staticWake[0] = (FrontendPlugin_dispatch_WRITE_RD_0 && FrontendPlugin_dispatch_LATENCY_0_0);
  assign DispatchPlugin_logic_pop_0_portEventFull = {DispatchPlugin_logic_queue_io_schedules_0_payload_event[7],{DispatchPlugin_logic_queue_io_schedules_0_payload_event[6],{DispatchPlugin_logic_queue_io_schedules_0_payload_event[5],{DispatchPlugin_logic_queue_io_schedules_0_payload_event[4],{DispatchPlugin_logic_queue_io_schedules_0_payload_event[3],{DispatchPlugin_logic_queue_io_schedules_0_payload_event[2],{DispatchPlugin_logic_queue_io_schedules_0_payload_event[1],DispatchPlugin_logic_queue_io_schedules_0_payload_event[0]}}}}}}};
  assign DispatchPlugin_logic_pop_0_stagesList_0_valid = DispatchPlugin_logic_queue_io_schedules_0_valid;
  assign DispatchPlugin_logic_pop_0_stagesList_0_OH = DispatchPlugin_logic_pop_0_portEventFull;
  assign DispatchPlugin_logic_pop_0_stagesList_0_OFFSET = DispatchPlugin_logic_ptr_current;
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT = DispatchPlugin_logic_pop_0_stagesList_0_OH[3];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_1 = DispatchPlugin_logic_pop_0_stagesList_0_OH[5];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_2 = DispatchPlugin_logic_pop_0_stagesList_0_OH[6];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3 = DispatchPlugin_logic_pop_0_stagesList_0_OH[7];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_4 = (((DispatchPlugin_logic_pop_0_stagesList_0_OH[1] || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3);
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_5 = (((DispatchPlugin_logic_pop_0_stagesList_0_OH[2] || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3);
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_6 = (((DispatchPlugin_logic_pop_0_stagesList_0_OH[4] || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3);
  assign DispatchPlugin_logic_pop_0_stagesList_0_UINT = {_zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_6,{_zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_5,_zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_4}};
  assign DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID = (_zz_DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID + DispatchPlugin_logic_pop_0_stagesList_1_OFFSET);
  assign DispatchPlugin_logic_pop_0_stagesList_0_LATENCY_0 = (|(DispatchPlugin_logic_pop_0_stagesList_0_OH & DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0));
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[1 : 0];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[3 : 2];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[5 : 4];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[7 : 6];
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0 = ((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0[0] ? DispatchPlugin_logic_queue_io_contexts_0_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0[1] ? DispatchPlugin_logic_queue_io_contexts_1_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1 = ((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1[0] ? DispatchPlugin_logic_queue_io_contexts_2_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1[1] ? DispatchPlugin_logic_queue_io_contexts_3_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2 = ((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2[0] ? DispatchPlugin_logic_queue_io_contexts_4_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2[1] ? DispatchPlugin_logic_queue_io_contexts_5_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3 = ((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3[0] ? DispatchPlugin_logic_queue_io_contexts_6_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3[1] ? DispatchPlugin_logic_queue_io_contexts_7_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_1_PHYS_RD = ((DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_0 | DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_1) | (DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_2 | DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_3));
  assign ALU0_ExecutionUnitBase_pipeline_push_port_valid = DispatchPlugin_logic_pop_0_stagesList_1_valid;
  assign ALU0_ExecutionUnitBase_pipeline_push_port_robId = DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_push_port_physRd = DispatchPlugin_logic_pop_0_stagesList_1_PHYS_RD;
  assign toplevel_DispatchPlugin_logic_queue_io_schedules_0_fire = (DispatchPlugin_logic_queue_io_schedules_0_valid && DispatchPlugin_logic_pop_0_stagesList_0_ready);
  assign DispatchPlugin_logic_pop_0_wake_L0_mask = (toplevel_DispatchPlugin_logic_queue_io_schedules_0_fire ? DispatchPlugin_logic_pop_0_portEventFull : 8'h00);
  assign DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid = (DispatchPlugin_logic_pop_0_stagesList_1_valid && DispatchPlugin_logic_pop_0_stagesList_1_LATENCY_0);
  assign DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical = DispatchPlugin_logic_pop_0_stagesList_1_PHYS_RD;
  assign DispatchPlugin_logic_pop_0_stagesList_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_0_stagesList_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_0_stagesList_0_ready = 1'b1;
  assign DispatchPlugin_logic_pop_1_portEventFull = {DispatchPlugin_logic_queue_io_schedules_1_payload_event[7],{DispatchPlugin_logic_queue_io_schedules_1_payload_event[6],{DispatchPlugin_logic_queue_io_schedules_1_payload_event[5],{DispatchPlugin_logic_queue_io_schedules_1_payload_event[4],{DispatchPlugin_logic_queue_io_schedules_1_payload_event[3],{DispatchPlugin_logic_queue_io_schedules_1_payload_event[2],{DispatchPlugin_logic_queue_io_schedules_1_payload_event[1],DispatchPlugin_logic_queue_io_schedules_1_payload_event[0]}}}}}}};
  assign DispatchPlugin_logic_pop_1_stagesList_0_valid = DispatchPlugin_logic_queue_io_schedules_1_valid;
  assign DispatchPlugin_logic_pop_1_stagesList_0_OH = DispatchPlugin_logic_pop_1_portEventFull;
  assign DispatchPlugin_logic_pop_1_stagesList_0_OFFSET = DispatchPlugin_logic_ptr_current;
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT = DispatchPlugin_logic_pop_1_stagesList_0_OH[3];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_1 = DispatchPlugin_logic_pop_1_stagesList_0_OH[5];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_2 = DispatchPlugin_logic_pop_1_stagesList_0_OH[6];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3 = DispatchPlugin_logic_pop_1_stagesList_0_OH[7];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_4 = (((DispatchPlugin_logic_pop_1_stagesList_0_OH[1] || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3);
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_5 = (((DispatchPlugin_logic_pop_1_stagesList_0_OH[2] || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3);
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_6 = (((DispatchPlugin_logic_pop_1_stagesList_0_OH[4] || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3);
  assign DispatchPlugin_logic_pop_1_stagesList_0_UINT = {_zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_6,{_zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_5,_zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_4}};
  assign DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID = (_zz_DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID + DispatchPlugin_logic_pop_1_stagesList_1_OFFSET);
  assign DispatchPlugin_logic_pop_1_stagesList_0_LATENCY_0 = (|(DispatchPlugin_logic_pop_1_stagesList_0_OH & DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0));
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_0 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[1 : 0];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_1 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[3 : 2];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_2 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[5 : 4];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_3 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[7 : 6];
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_0 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_0[0] ? DispatchPlugin_logic_queue_io_contexts_0_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_0[1] ? DispatchPlugin_logic_queue_io_contexts_1_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_1 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_1[0] ? DispatchPlugin_logic_queue_io_contexts_2_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_1[1] ? DispatchPlugin_logic_queue_io_contexts_3_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_2 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_2[0] ? DispatchPlugin_logic_queue_io_contexts_4_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_2[1] ? DispatchPlugin_logic_queue_io_contexts_5_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_3 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_3[0] ? DispatchPlugin_logic_queue_io_contexts_6_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_3[1] ? DispatchPlugin_logic_queue_io_contexts_7_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RD = ((DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_0 | DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_1) | (DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_2 | DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_3));
  assign EU0_ExecutionUnitBase_pipeline_push_port_valid = DispatchPlugin_logic_pop_1_stagesList_1_valid;
  assign EU0_ExecutionUnitBase_pipeline_push_port_robId = DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_push_port_physRd = DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RD;
  assign DispatchPlugin_logic_pop_1_stagesList_1_haltRequest_DispatchPlugin_l292 = (! EU0_ExecutionUnitBase_pipeline_push_port_ready);
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_0 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[1 : 0];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_1 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[3 : 2];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_2 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[5 : 4];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_3 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[7 : 6];
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_0 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_0[0] ? DispatchPlugin_logic_queue_io_contexts_0_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_0[1] ? DispatchPlugin_logic_queue_io_contexts_1_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_1 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_1[0] ? DispatchPlugin_logic_queue_io_contexts_2_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_1[1] ? DispatchPlugin_logic_queue_io_contexts_3_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_2 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_2[0] ? DispatchPlugin_logic_queue_io_contexts_4_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_2[1] ? DispatchPlugin_logic_queue_io_contexts_5_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_3 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_3[0] ? DispatchPlugin_logic_queue_io_contexts_6_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_3[1] ? DispatchPlugin_logic_queue_io_contexts_7_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RS_0 = ((DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_0 | DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_1) | (DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_2 | DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_3));
  assign EU0_ExecutionUnitBase_pipeline_push_port_context_0 = DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RS_0;
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_0 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[1 : 0];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_1 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[3 : 2];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_2 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[5 : 4];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_3 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[7 : 6];
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_0 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_0[0] ? DispatchPlugin_logic_queue_io_contexts_0_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_0[1] ? DispatchPlugin_logic_queue_io_contexts_1_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_1 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_1[0] ? DispatchPlugin_logic_queue_io_contexts_2_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_1[1] ? DispatchPlugin_logic_queue_io_contexts_3_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_2 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_2[0] ? DispatchPlugin_logic_queue_io_contexts_4_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_2[1] ? DispatchPlugin_logic_queue_io_contexts_5_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_3 = ((_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_3[0] ? DispatchPlugin_logic_queue_io_contexts_6_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_3[1] ? DispatchPlugin_logic_queue_io_contexts_7_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RS_1 = ((DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_0 | DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_1) | (DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_2 | DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_3));
  assign EU0_ExecutionUnitBase_pipeline_push_port_context_1 = DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RS_1;
  assign DispatchPlugin_logic_pop_1_stagesList_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_1_stagesList_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_1_stagesList_0_ready = DispatchPlugin_logic_pop_1_stagesList_0_ready_output;
  always @(*) begin
    DispatchPlugin_logic_pop_1_stagesList_1_ready = 1'b1;
    if(when_Pipeline_l278_5) begin
      DispatchPlugin_logic_pop_1_stagesList_1_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_5 = (|DispatchPlugin_logic_pop_1_stagesList_1_haltRequest_DispatchPlugin_l292);
  always @(*) begin
    DispatchPlugin_logic_pop_1_stagesList_0_ready_output = DispatchPlugin_logic_pop_1_stagesList_1_ready;
    if(when_Connection_l74_4) begin
      DispatchPlugin_logic_pop_1_stagesList_0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_4 = (! DispatchPlugin_logic_pop_1_stagesList_1_valid);
  assign DispatchPlugin_logic_wake_dynamic_offseted_0_valid = Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_valid;
  assign DispatchPlugin_logic_wake_dynamic_offseted_0_payload = _zz_DispatchPlugin_logic_wake_dynamic_offseted_0_payload[2:0];
  assign DispatchPlugin_logic_wake_dynamic_offseted_1_valid = Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_valid;
  assign DispatchPlugin_logic_wake_dynamic_offseted_1_payload = _zz_DispatchPlugin_logic_wake_dynamic_offseted_1_payload[2:0];
  assign DispatchPlugin_logic_wake_dynamic_offseted_2_valid = Lsu2Plugin_logic_special_wakeRob_valid;
  assign DispatchPlugin_logic_wake_dynamic_offseted_2_payload = _zz_DispatchPlugin_logic_wake_dynamic_offseted_2_payload[2:0];
  assign DispatchPlugin_logic_wake_dynamic_offseted_3_valid = EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_valid;
  assign DispatchPlugin_logic_wake_dynamic_offseted_3_payload = _zz_DispatchPlugin_logic_wake_dynamic_offseted_3_payload[2:0];
  assign DispatchPlugin_logic_wake_dynamic_masks_0 = ((DispatchPlugin_logic_wake_dynamic_offseted_0_valid ? 8'hff : 8'h00) & _zz_DispatchPlugin_logic_wake_dynamic_masks_0);
  assign DispatchPlugin_logic_wake_dynamic_masks_1 = ((DispatchPlugin_logic_wake_dynamic_offseted_1_valid ? 8'hff : 8'h00) & _zz_DispatchPlugin_logic_wake_dynamic_masks_1);
  assign DispatchPlugin_logic_wake_dynamic_masks_2 = ((DispatchPlugin_logic_wake_dynamic_offseted_2_valid ? 8'hff : 8'h00) & _zz_DispatchPlugin_logic_wake_dynamic_masks_2);
  assign DispatchPlugin_logic_wake_dynamic_masks_3 = ((DispatchPlugin_logic_wake_dynamic_offseted_3_valid ? 8'hff : 8'h00) & _zz_DispatchPlugin_logic_wake_dynamic_masks_3);
  assign DispatchPlugin_logic_wake_statics_0_popMask = (DispatchPlugin_logic_pop_0_wake_L0_mask & DispatchPlugin_logic_queueStaticWakeTransposed_0);
  assign DispatchPlugin_logic_wake_statics_0_history_0 = DispatchPlugin_logic_wake_statics_0_popMask;
  assign DispatchPlugin_logic_wake_optReduce_relaxed = ((DispatchPlugin_logic_wake_dynamic_masks_0 | DispatchPlugin_logic_wake_dynamic_masks_1) | (DispatchPlugin_logic_wake_dynamic_masks_2 | DispatchPlugin_logic_wake_dynamic_masks_3));
  assign DispatchPlugin_logic_wake_optReduce_reduced = (DispatchPlugin_logic_wake_optReduce_relaxed | DispatchPlugin_logic_wake_statics_0_history_0);
  assign DispatchPlugin_logic_whitebox_issuePorts_0_valid = (ALU0_ExecutionUnitBase_pipeline_push_port_valid && 1'b1);
  assign DispatchPlugin_logic_whitebox_issuePorts_0_payload_robId = ALU0_ExecutionUnitBase_pipeline_push_port_robId;
  assign DispatchPlugin_logic_whitebox_issuePorts_0_payload_physRd = ALU0_ExecutionUnitBase_pipeline_push_port_physRd;
  assign DispatchPlugin_logic_whitebox_issuePorts_1_valid = (EU0_ExecutionUnitBase_pipeline_push_port_valid && EU0_ExecutionUnitBase_pipeline_push_port_ready);
  assign DispatchPlugin_logic_whitebox_issuePorts_1_payload_robId = EU0_ExecutionUnitBase_pipeline_push_port_robId;
  assign DispatchPlugin_logic_whitebox_issuePorts_1_payload_physRd = EU0_ExecutionUnitBase_pipeline_push_port_physRd;
  assign DispatchPlugin_logic_whitebox_issuePorts_1_payload_context_0 = EU0_ExecutionUnitBase_pipeline_push_port_context_0;
  assign DispatchPlugin_logic_whitebox_issuePorts_1_payload_context_1 = EU0_ExecutionUnitBase_pipeline_push_port_context_1;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_valid = (|{EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid,Lsu2Plugin_setup_regfilePorts_0_write_valid});
  assign _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0 = {EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid,Lsu2Plugin_setup_regfilePorts_0_write_valid};
  assign _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_1 = _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0[0];
  always @(*) begin
    _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_2[0] = (_zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_1 && (! 1'b0));
    _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_2[1] = (_zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0[1] && (! _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_1));
  end

  assign _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_3 = _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_2;
  assign integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0 = _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_3[0];
  assign integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_1 = _zz_integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0_3[1];
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_address = ((integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0 ? Lsu2Plugin_setup_regfilePorts_0_write_address : 6'h00) | (integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_1 ? EU0_ExecutionUnitBase_pipeline_writeBack_0_write_address : 6'h00));
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_data = ((integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0 ? Lsu2Plugin_setup_regfilePorts_0_write_data : 32'h00000000) | (integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_1 ? EU0_ExecutionUnitBase_pipeline_writeBack_0_write_data : 32'h00000000));
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_robId = ((integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_0 ? Lsu2Plugin_setup_regfilePorts_0_write_robId : 4'b0000) | (integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_1 ? EU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId : 4'b0000));
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_ready = integer_RegFilePlugin_logic_writeMerges_0_multiple_oh_1;
  assign integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid = Lsu2Plugin_setup_regfilePorts_0_write_valid;
  assign integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address = Lsu2Plugin_setup_regfilePorts_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data = Lsu2Plugin_setup_regfilePorts_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_valid = (|ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid);
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_address = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_data = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_robId = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  assign integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid;
  assign integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  always @(*) begin
    ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = integer_RegFilePlugin_logic_regfile_latches_io_reads_0_data;
    if(when_RegFilePlugin_l327) begin
      ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = (_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data ? integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data : integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data);
    end
  end

  always @(*) begin
    ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = integer_RegFilePlugin_logic_regfile_latches_io_reads_1_data;
    if(when_RegFilePlugin_l327_1) begin
      ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = (_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data ? integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data : integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data);
    end
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = integer_RegFilePlugin_logic_regfile_latches_io_reads_2_data;
    if(when_RegFilePlugin_l327_2) begin
      EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = (_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data ? integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data : integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data);
    end
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = integer_RegFilePlugin_logic_regfile_latches_io_reads_3_data;
    if(when_RegFilePlugin_l327_3) begin
      EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = (_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data ? integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data : integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data);
    end
  end

  assign _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address));
  assign when_RegFilePlugin_l327 = (|{(integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address)),_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data});
  assign _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address));
  assign when_RegFilePlugin_l327_1 = (|{(integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address)),_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data});
  assign _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address));
  assign when_RegFilePlugin_l327_2 = (|{(integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address)),_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data});
  assign _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address));
  assign when_RegFilePlugin_l327_3 = (|{(integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address)),_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data});
  assign integer_write_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  assign integer_write_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  assign integer_write_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  assign integer_write_0_robId = integer_RegFilePlugin_logic_writeMerges_0_bus_robId;
  assign integer_write_1_valid = integer_RegFilePlugin_logic_writeMerges_1_bus_valid;
  assign integer_write_1_address = integer_RegFilePlugin_logic_writeMerges_1_bus_address;
  assign integer_write_1_data = integer_RegFilePlugin_logic_writeMerges_1_bus_data;
  assign integer_write_1_robId = integer_RegFilePlugin_logic_writeMerges_1_bus_robId;
  assign AguPlugin_setup_port_payload_earlySample = EU0_ExecutionUnitBase_pipeline_fetch_0_ready;
  assign AguPlugin_setup_port_payload_earlyPc = EU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  assign RobPlugin_logic_completionMem_targetWrite_valid = FrontendPlugin_allocated_isFireing;
  assign RobPlugin_logic_completionMem_targetWrite_payload_address = FrontendPlugin_allocated_ROB_ID;
  assign RobPlugin_logic_completionMem_init_0_robId = FrontendPlugin_allocated_ROB_ID;
  assign RobPlugin_logic_completionMem_targetWrite_payload_data[0] = (^{RobPlugin_logic_completionMem_hits_3_spinal_port0[0],{RobPlugin_logic_completionMem_hits_2_spinal_port0[0],{RobPlugin_logic_completionMem_hits_1_spinal_port0[0],RobPlugin_logic_completionMem_hits_0_spinal_port0[0]}}});
  assign RobPlugin_logic_completionMem_reads_0_targetRead_data = RobPlugin_logic_completionMem_target_spinal_port1;
  assign RobPlugin_logic_completionMem_reads_0_targetRead_address = CommitPlugin_setup_robLineMask_line;
  assign _zz_CommitPlugin_setup_robLineMask_mask = CommitPlugin_setup_robLineMask_line;
  always @(*) begin
    CommitPlugin_setup_robLineMask_mask[0] = ((^{RobPlugin_logic_completionMem_hits_3_spinal_port3[0],{RobPlugin_logic_completionMem_hits_2_spinal_port3[0],{RobPlugin_logic_completionMem_hits_1_spinal_port3[0],RobPlugin_logic_completionMem_hits_0_spinal_port3[0]}}}) != RobPlugin_logic_completionMem_reads_0_targetRead_data[0]);
    if(when_RobPlugin_l118) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_1) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_2) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_3) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l123) begin
      CommitPlugin_setup_robLineMask_mask = 1'b0;
    end
  end

  assign _zz_when_RobPlugin_l118 = CommitPlugin_setup_robLineMask_line;
  assign when_RobPlugin_l118 = (Lsu2Plugin_setup_sharedCompletion_valid && (Lsu2Plugin_setup_sharedCompletion_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_1 = (Lsu2Plugin_setup_specialCompletion_valid && (Lsu2Plugin_setup_specialCompletion_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_2 = (ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid && (ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_3 = (EU0_ExecutionUnitBase_pipeline_completion_0_port_valid && (EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l123 = (FrontendPlugin_allocated_isFireing && (FrontendPlugin_allocated_ROB_ID == CommitPlugin_setup_robLineMask_line));
  assign _zz_CommitPlugin_logic_commit_active = CommitPlugin_logic_ptr_commit[3 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_mask_0 = CommitPlugin_logic_free_port_payload_robId;
  assign integer_RfAllocationPlugin_logic_push_mask_0 = _zz_integer_RfAllocationPlugin_logic_push_mask_0_1[0];
  assign _zz_commit_pc_0 = CommitPlugin_logic_commit_event_robId;
  assign _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc = CommitPlugin_logic_commit_reschedulePort_payload_robId;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC = ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0 = CommitPlugin_logic_commit_event_robId;
  assign integer_RfTranslationPlugin_logic_onCommit_writeRd_0 = _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1[0];
  assign _zz_integer_RfAllocationPlugin_logic_push_writeRd_0 = CommitPlugin_logic_free_port_payload_robId;
  assign integer_RfAllocationPlugin_logic_push_writeRd_0 = _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0 = CommitPlugin_logic_commit_event_robId;
  assign integer_RfTranslationPlugin_logic_onCommit_physRd_0 = _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_1[5 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0 = CommitPlugin_logic_free_port_payload_robId;
  assign integer_RfAllocationPlugin_logic_push_physicalRdNew_0 = _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_1[5 : 0];
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0 = CommitPlugin_logic_commit_event_robId;
  assign integer_RfTranslationPlugin_logic_onCommit_archRd_0 = _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_1[4 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0 = CommitPlugin_logic_free_port_payload_robId;
  assign integer_RfAllocationPlugin_logic_push_physicalRdOld_0 = _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_1[5 : 0];
  assign _zz_BranchContextPlugin_logic_onCommit_isBranch_0 = CommitPlugin_logic_commit_event_robId;
  assign BranchContextPlugin_logic_onCommit_isBranch_0 = _zz_BranchContextPlugin_logic_onCommit_isBranch_0_1[0];
  assign _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0 = CommitPlugin_logic_commit_event_robId;
  assign HistoryPlugin_logic_onCommit_isConditionalBranch_0 = _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1[0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch = CommitPlugin_logic_reschedule_reschedulePort_payload_robId;
  assign _zz_HistoryPlugin_logic_onCommit_isTaken_0 = CommitPlugin_logic_commit_event_robId;
  assign HistoryPlugin_logic_onCommit_isTaken_0 = _zz_HistoryPlugin_logic_onCommit_isTaken_0_1[0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken = CommitPlugin_logic_reschedule_reschedulePort_payload_robId;
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory = CommitPlugin_logic_reschedule_reschedulePort_payload_robId;
  assign _zz_DecoderPredictionPlugin_logic_ras_healPush = CommitPlugin_logic_reschedule_reschedulePort_payload_robId;
  assign _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0 = CommitPlugin_logic_commit_event_robId;
  assign Lsu2Plugin_logic_lq_onCommit_lqAlloc_0 = _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_1[0];
  assign _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0 = CommitPlugin_logic_commit_event_robId;
  assign Lsu2Plugin_logic_sq_onCommit_sqAlloc_0 = _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0 = ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1 = ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  assign RobPlugin_logic_whitebox_completionsPorts_0_valid = Lsu2Plugin_setup_sharedCompletion_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_0_payload_id = Lsu2Plugin_setup_sharedCompletion_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_1_valid = Lsu2Plugin_setup_specialCompletion_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_1_payload_id = Lsu2Plugin_setup_specialCompletion_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_2_valid = ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_2_payload_id = ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_3_valid = EU0_ExecutionUnitBase_pipeline_completion_0_port_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_3_payload_id = EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_valid = (((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_WRITE_RD_0) && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_payload_robId = (FrontendPlugin_dispatch_ROB_ID | 4'b0000);
  always @(*) begin
    RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_valid = (DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid && 1'b1);
    if(RfDependencyPlugin_logic_forRf_integer_init_busy) begin
      RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_valid = 1'b1;
    end
  end

  always @(*) begin
    RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_payload_physical = DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical;
    if(RfDependencyPlugin_logic_forRf_integer_init_busy) begin
      RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_payload_physical = RfDependencyPlugin_logic_forRf_integer_init_counter[5:0];
    end
  end

  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_1_valid = (Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_2_valid = (Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_3_valid = (Lsu2Plugin_logic_special_wakeRf_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_4_valid = (EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_init_busy = (! RfDependencyPlugin_logic_forRf_integer_init_counter[6]);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_cmd_valid = ((FrontendPlugin_dispatch_valid && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && FrontendPlugin_dispatch_READ_RS_0_0);
  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = 1'bx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_enable;
  end

  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0 = 4'bxxxx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_rob;
  end

  always @(*) begin
    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0;
    if(when_RfDependencyPlugin_l228) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = 1'b0;
    end
    if(when_RfDependencyPlugin_l232) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = 1'b0;
    end
  end

  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0;
  assign when_RfDependencyPlugin_l228 = ((DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_0_0)) && 1'b1);
  assign when_RfDependencyPlugin_l232 = (! FrontendPlugin_dispatch_READ_RS_0_0);
  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_0 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 && (! FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_0));
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_cmd_valid = ((FrontendPlugin_dispatch_valid && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && FrontendPlugin_dispatch_READ_RS_1_0);
  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = 1'bx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_enable;
  end

  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0 = 4'bxxxx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_rob;
  end

  always @(*) begin
    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0;
    if(when_RfDependencyPlugin_l228_1) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = 1'b0;
    end
    if(when_RfDependencyPlugin_l232_1) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = 1'b0;
    end
  end

  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0;
  assign when_RfDependencyPlugin_l228_1 = ((DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_1_0)) && 1'b1);
  assign when_RfDependencyPlugin_l232_1 = (! FrontendPlugin_dispatch_READ_RS_1_0);
  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_0 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 && (! FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_0));
  assign FrontendPlugin_isBusy = (|{FrontendPlugin_dispatch_valid,{FrontendPlugin_allocated_valid,{FrontendPlugin_serialized_valid,{FrontendPlugin_decoded_valid,FrontendPlugin_decompressed_valid}}}});
  assign FrontendPlugin_isBusyAfterDecode = (|{FrontendPlugin_dispatch_valid,{FrontendPlugin_allocated_valid,FrontendPlugin_serialized_valid}});
  assign FrontendPlugin_dispatch_isFlushed = CommitPlugin_logic_reschedule_reschedulePort_valid;
  assign FrontendPlugin_allocated_isFlushed = CommitPlugin_logic_reschedule_reschedulePort_valid;
  assign when_Connection_l66 = (|{CommitPlugin_logic_reschedule_reschedulePort_valid,(DecoderPredictionPlugin_setup_decodeJump_valid && FrontendPlugin_serialized_ready)});
  assign FrontendPlugin_serialized_isFlushed = when_Connection_l66;
  assign _zz_FrontendPlugin_decompressed_isFlushed = (|{when_Connection_l66,_zz_FrontendPlugin_decoded_isFlushingRoot});
  assign FrontendPlugin_decoded_isFlushed = _zz_FrontendPlugin_decompressed_isFlushed;
  assign FrontendPlugin_decompressed_isFlushed = _zz_FrontendPlugin_decompressed_isFlushed;
  assign FrontendPlugin_aligned_isFlushed = _zz_FrontendPlugin_decompressed_isFlushed;
  assign FrontendPlugin_decoded_isFlushingRoot = (|_zz_FrontendPlugin_decoded_isFlushingRoot);
  assign FrontendPlugin_dispatch_isFlushingRoot = (|CommitPlugin_logic_reschedule_reschedulePort_valid);
  assign FrontendPlugin_aligned_ready = FrontendPlugin_aligned_ready_output;
  assign FrontendPlugin_decompressed_ready = FrontendPlugin_decompressed_ready_output;
  always @(*) begin
    _zz_FrontendPlugin_serialized_valid = FrontendPlugin_decoded_valid;
    if(FrontendPlugin_decoded_isFlushingRoot) begin
      _zz_FrontendPlugin_serialized_valid = 1'b0;
    end
    if(when_Pipeline_l278_6) begin
      _zz_FrontendPlugin_serialized_valid = 1'b0;
    end
  end

  always @(*) begin
    FrontendPlugin_decoded_ready = FrontendPlugin_decoded_ready_output;
    if(when_Pipeline_l278_6) begin
      FrontendPlugin_decoded_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_6 = (|{FrontendPlugin_decoded_haltRequest_DecoderPlugin_l325,FrontendPlugin_decoded_haltRequest_DecoderPlugin_l324});
  assign FrontendPlugin_serialized_ready = FrontendPlugin_serialized_ready_output;
  always @(*) begin
    _zz_FrontendPlugin_dispatch_valid = FrontendPlugin_allocated_valid;
    if(when_Pipeline_l278_7) begin
      _zz_FrontendPlugin_dispatch_valid = 1'b0;
    end
  end

  always @(*) begin
    FrontendPlugin_allocated_ready = FrontendPlugin_allocated_ready_output;
    if(when_Pipeline_l278_7) begin
      FrontendPlugin_allocated_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_7 = (|{FrontendPlugin_allocated_haltRequest_FrontendPlugin_l67,{FrontendPlugin_allocated_haltRequest_CommitPlugin_l95,{FrontendPlugin_allocated_haltRequest_BranchContextPlugin_l111,FrontendPlugin_allocated_haltRequest_RfAllocationPlugin_l55}}});
  always @(*) begin
    FrontendPlugin_dispatch_ready = 1'b1;
    if(when_Pipeline_l278_8) begin
      FrontendPlugin_dispatch_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_8 = (|{FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l196,{FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l195,{FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l187,{FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l1838,FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l620}}}});
  assign FrontendPlugin_serialized_ready_output = FrontendPlugin_allocated_ready;
  assign FrontendPlugin_allocated_valid = FrontendPlugin_serialized_valid;
  assign FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_0 = FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0;
  assign FrontendPlugin_allocated_Frontend_MICRO_OP_0 = FrontendPlugin_serialized_Frontend_MICRO_OP_0;
  assign FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_0 = FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0;
  assign FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_0 = FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0;
  assign FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_0 = FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0;
  assign FrontendPlugin_allocated_BRANCH_SEL_0 = FrontendPlugin_serialized_BRANCH_SEL_0;
  assign FrontendPlugin_allocated_BRANCH_EARLY_0_taken = FrontendPlugin_serialized_BRANCH_EARLY_0_taken;
  assign FrontendPlugin_allocated_BRANCH_EARLY_0_pc = FrontendPlugin_serialized_BRANCH_EARLY_0_pc;
  assign FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0 = FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0;
  assign FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_0 = FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_0;
  assign FrontendPlugin_allocated_Prediction_IS_BRANCH_0 = FrontendPlugin_serialized_Prediction_IS_BRANCH_0;
  assign FrontendPlugin_allocated_FETCH_ID_0 = FrontendPlugin_serialized_FETCH_ID_0;
  assign FrontendPlugin_allocated_WRITE_RD_0 = FrontendPlugin_serialized_WRITE_RD_0;
  assign FrontendPlugin_allocated_PC_0 = FrontendPlugin_serialized_PC_0;
  assign FrontendPlugin_allocated_ARCH_RD_0 = FrontendPlugin_serialized_ARCH_RD_0;
  assign FrontendPlugin_allocated_ARCH_RS_0_0 = FrontendPlugin_serialized_ARCH_RS_0_0;
  assign FrontendPlugin_allocated_READ_RS_0_0 = FrontendPlugin_serialized_READ_RS_0_0;
  assign FrontendPlugin_allocated_ARCH_RS_1_0 = FrontendPlugin_serialized_ARCH_RS_1_0;
  assign FrontendPlugin_allocated_READ_RS_1_0 = FrontendPlugin_serialized_READ_RS_1_0;
  assign FrontendPlugin_allocated_BRANCH_HISTORY_0 = FrontendPlugin_serialized_BRANCH_HISTORY_0;
  assign FrontendPlugin_allocated_OP_ID = FrontendPlugin_serialized_OP_ID;
  assign FrontendPlugin_allocated_LQ_ALLOC_0 = FrontendPlugin_serialized_LQ_ALLOC_0;
  assign FrontendPlugin_allocated_SQ_ALLOC_0 = FrontendPlugin_serialized_SQ_ALLOC_0;
  assign FrontendPlugin_allocated_GSHARE_COUNTER_0_0 = FrontendPlugin_serialized_GSHARE_COUNTER_0_0;
  assign FrontendPlugin_allocated_ALU0_SEL_0 = FrontendPlugin_serialized_ALU0_SEL_0;
  assign FrontendPlugin_allocated_EU0_SEL_0 = FrontendPlugin_serialized_EU0_SEL_0;
  always @(*) begin
    FrontendPlugin_allocated_ready_output = FrontendPlugin_dispatch_ready;
    if(when_Connection_l74_5) begin
      FrontendPlugin_allocated_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_5 = (! FrontendPlugin_dispatch_valid);
  assign FrontendPlugin_aligned_ready_output = FrontendPlugin_decompressed_ready;
  assign FrontendPlugin_decompressed_valid = FrontendPlugin_aligned_valid;
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_0 = FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_0;
  assign FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_0 = FrontendPlugin_aligned_Frontend_MASK_ALIGNED_0;
  assign FrontendPlugin_decompressed_PC_0 = FrontendPlugin_aligned_PC_0;
  assign FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_0 = FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0;
  assign FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_0 = FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  assign FrontendPlugin_decompressed_BRANCH_HISTORY_0 = FrontendPlugin_aligned_BRANCH_HISTORY_0;
  assign FrontendPlugin_decompressed_GSHARE_COUNTER_0_0 = FrontendPlugin_aligned_GSHARE_COUNTER_0_0;
  assign FrontendPlugin_decompressed_FETCH_ID_0 = FrontendPlugin_aligned_FETCH_ID_0;
  assign FrontendPlugin_decompressed_Frontend_FETCH_FAULT_0 = FrontendPlugin_aligned_Frontend_FETCH_FAULT_0;
  assign FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_0 = FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0;
  assign FrontendPlugin_decompressed_ready_output = FrontendPlugin_decoded_ready;
  assign FrontendPlugin_decoded_valid = FrontendPlugin_decompressed_valid;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_0;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_0 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_0;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_0 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_0;
  assign FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_0 = FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_0;
  assign FrontendPlugin_decoded_GSHARE_COUNTER_0_0 = FrontendPlugin_decompressed_GSHARE_COUNTER_0_0;
  assign FrontendPlugin_decoded_FETCH_ID_0 = FrontendPlugin_decompressed_FETCH_ID_0;
  assign FrontendPlugin_decoded_Frontend_MASK_ALIGNED_0 = FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_0;
  assign FrontendPlugin_decoded_Frontend_FETCH_FAULT_0 = FrontendPlugin_decompressed_Frontend_FETCH_FAULT_0;
  assign FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_0 = FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_0;
  assign FrontendPlugin_decoded_PC_0 = FrontendPlugin_decompressed_PC_0;
  assign FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_0 = FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  assign FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_0 = FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_0;
  assign FrontendPlugin_decoded_BRANCH_HISTORY_0 = FrontendPlugin_decompressed_BRANCH_HISTORY_0;
  always @(*) begin
    FrontendPlugin_decoded_ready_output = FrontendPlugin_serialized_ready;
    if(when_Connection_l74_6) begin
      FrontendPlugin_decoded_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_6 = (! FrontendPlugin_serialized_valid);
  assign PcPlugin_logic_init_booted = PcPlugin_logic_init_counter[6];
  always @(*) begin
    PcPlugin_logic_fetchPc_correction = 1'b0;
    if(PcPlugin_logic_jump_pcLoad_valid) begin
      PcPlugin_logic_fetchPc_correction = 1'b1;
    end
  end

  assign PcPlugin_logic_fetchPc_output_fire = (PcPlugin_logic_fetchPc_output_valid && PcPlugin_logic_fetchPc_output_ready);
  assign PcPlugin_logic_fetchPc_corrected = (PcPlugin_logic_fetchPc_correction || PcPlugin_logic_fetchPc_correctionReg);
  assign PcPlugin_logic_fetchPc_pcRegPropagate = 1'b0;
  assign when_PcPlugin_l84 = (PcPlugin_logic_fetchPc_correction || PcPlugin_logic_fetchPc_pcRegPropagate);
  assign when_PcPlugin_l84_1 = ((! PcPlugin_logic_fetchPc_output_valid) && PcPlugin_logic_fetchPc_output_ready);
  always @(*) begin
    PcPlugin_logic_fetchPc_pc = (PcPlugin_logic_fetchPc_pcReg + _zz_PcPlugin_logic_fetchPc_pc);
    if(PcPlugin_logic_jump_pcLoad_valid) begin
      PcPlugin_logic_fetchPc_pc = PcPlugin_logic_jump_pcLoad_payload_pc;
    end
    PcPlugin_logic_fetchPc_pc[0] = 1'b0;
    PcPlugin_logic_fetchPc_pc[1] = 1'b0;
  end

  always @(*) begin
    PcPlugin_logic_fetchPc_flushed = 1'b0;
    if(PcPlugin_logic_jump_pcLoad_valid) begin
      PcPlugin_logic_fetchPc_flushed = 1'b1;
    end
  end

  assign when_PcPlugin_l100 = (PcPlugin_logic_init_booted && ((PcPlugin_logic_fetchPc_output_ready || PcPlugin_logic_fetchPc_correction) || PcPlugin_logic_fetchPc_pcRegPropagate));
  assign PcPlugin_logic_fetchPc_fetcherHalt = 1'b0;
  assign PcPlugin_logic_fetchPc_output_valid = ((! PcPlugin_logic_fetchPc_fetcherHalt) && PcPlugin_logic_init_booted);
  assign PcPlugin_logic_fetchPc_output_payload = PcPlugin_logic_fetchPc_pc;
  assign PcPlugin_logic_fetchPc_output_ready = FetchPlugin_stages_0_ready;
  assign FetchPlugin_stages_0_valid = PcPlugin_logic_fetchPc_output_valid;
  assign FetchPlugin_stages_0_Fetch_FETCH_PC = PcPlugin_logic_fetchPc_output_payload;
  always @(*) begin
    FetchPlugin_stages_1_Fetch_FETCH_PC_INC = (FetchPlugin_stages_1_Fetch_FETCH_PC + 32'h00000004);
    FetchPlugin_stages_1_Fetch_FETCH_PC_INC[1 : 0] = 2'b00;
  end

  assign fetchLastFire = FetchPlugin_stages_2_isFireing;
  assign fetchLastId = FetchPlugin_stages_2_FETCH_ID;
  assign AlignerPlugin_setup_s2m_isFlushed = FrontendPlugin_aligned_isFlushed;
  assign when_Connection_l66_1 = (|{FrontendPlugin_aligned_isFlushed,_zz_FetchPlugin_stages_2_isFlushingRoot});
  assign FetchPlugin_stages_2_isFlushed = when_Connection_l66_1;
  assign FetchPlugin_stages_1_isRemoved = (FetchPlugin_stages_1_isFlushed || FetchPlugin_stages_1_isThrown);
  assign when_Connection_l54 = (|{when_Connection_l66_1,_zz_FetchPlugin_stages_1_isFlushingRoot});
  assign FetchPlugin_stages_1_isFlushed = when_Connection_l54;
  assign FetchPlugin_stages_1_isFlushingNext = BtbPlugin_logic_applyIt_doIt;
  assign FetchPlugin_stages_1_isThrown = 1'b0;
  assign FetchPlugin_stages_0_isFlushed = (when_Connection_l54 || (BtbPlugin_logic_applyIt_doIt && 1'b1));
  assign FetchPlugin_stages_1_isFlushingRoot = (|_zz_FetchPlugin_stages_1_isFlushingRoot);
  assign FetchPlugin_stages_2_isFlushingRoot = (|_zz_FetchPlugin_stages_2_isFlushingRoot);
  assign AlignerPlugin_setup_s2m_isFlushingRoot = 1'b0;
  always @(*) begin
    _zz_FetchPlugin_stages_1_valid = FetchPlugin_stages_0_valid;
    if(when_Pipeline_l278_9) begin
      _zz_FetchPlugin_stages_1_valid = 1'b0;
    end
  end

  always @(*) begin
    FetchPlugin_stages_0_ready = FetchPlugin_stages_0_ready_output;
    if(when_Pipeline_l278_9) begin
      FetchPlugin_stages_0_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_9 = (|{FetchPlugin_stages_0_haltRequest_MmuPlugin_l533,{FetchPlugin_stages_0_haltRequest_EnvCallPlugin_l138,{FetchPlugin_stages_0_haltRequest_PrivilegedPlugin_l975,{FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548,{FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l583,{FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552,{FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l476,FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l389}}}}}}});
  always @(*) begin
    _zz_FetchPlugin_stages_2_valid = FetchPlugin_stages_1_valid;
    if(FetchPlugin_stages_1_isFlushingRoot) begin
      _zz_FetchPlugin_stages_2_valid = 1'b0;
    end
  end

  assign FetchPlugin_stages_1_ready = FetchPlugin_stages_1_ready_output;
  always @(*) begin
    _zz_AlignerPlugin_setup_s2m_valid = FetchPlugin_stages_2_valid;
    if(FetchPlugin_stages_2_isFlushingRoot) begin
      _zz_AlignerPlugin_setup_s2m_valid = 1'b0;
    end
  end

  assign FetchPlugin_stages_2_ready = FetchPlugin_stages_2_ready_output;
  always @(*) begin
    AlignerPlugin_setup_s2m_ready = 1'b1;
    if(when_Pipeline_l278_10) begin
      AlignerPlugin_setup_s2m_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_10 = (|AlignerPlugin_setup_s2m_haltRequest_AlignerPlugin_l270);
  always @(*) begin
    FetchPlugin_stages_0_ready_output = FetchPlugin_stages_1_ready;
    if(when_Connection_l74_7) begin
      FetchPlugin_stages_0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_7 = (! FetchPlugin_stages_1_valid);
  always @(*) begin
    FetchPlugin_stages_1_ready_output = FetchPlugin_stages_2_ready;
    if(when_Connection_l74_8) begin
      FetchPlugin_stages_1_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_8 = (! FetchPlugin_stages_2_valid);
  assign FetchPlugin_stages_2_ready_output = (! FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid);
  assign AlignerPlugin_setup_s2m_valid = (_zz_AlignerPlugin_setup_s2m_valid || FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid);
  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_WORD = FetchPlugin_stages_2_Fetch_WORD_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_WORD = FetchPlugin_stages_2_Fetch_WORD;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_FETCH_PC = FetchPlugin_stages_2_Fetch_FETCH_PC_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_FETCH_PC = FetchPlugin_stages_2_Fetch_FETCH_PC;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_WORD_FAULT = FetchPlugin_stages_2_Fetch_WORD_FAULT_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_WORD_FAULT = FetchPlugin_stages_2_Fetch_WORD_FAULT;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE = FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE = FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_BRANCH_HISTORY = FetchPlugin_stages_2_BRANCH_HISTORY_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_BRANCH_HISTORY = FetchPlugin_stages_2_BRANCH_HISTORY;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_FETCH_ID = FetchPlugin_stages_2_FETCH_ID_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_FETCH_ID = FetchPlugin_stages_2_FETCH_ID;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID = FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID = FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_MASK_FRONT = FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_MASK_FRONT = FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT = FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT = FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_GSHARE_COUNTER_0 = FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_0;
    end else begin
      AlignerPlugin_setup_s2m_GSHARE_COUNTER_0 = FetchPlugin_stages_2_GSHARE_COUNTER_0;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_FETCH_PC_INC = FetchPlugin_stages_2_Fetch_FETCH_PC_INC_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_FETCH_PC_INC = FetchPlugin_stages_2_Fetch_FETCH_PC_INC;
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_stateReg;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
        if(PrivilegedPlugin_logic_rescheduleUnbuffered_valid) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_SETUP;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
        if(when_PrivilegedPlugin_l773) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ;
        end else begin
          case(PrivilegedPlugin_logic_reschedule_payload_cause)
            4'b1001 : begin
              PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC;
            end
            4'b1010 : begin
              PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC;
            end
            4'b1000 : begin
              PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_EPC_READ;
            end
            default : begin
              PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ;
            end
          endcase
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        if(PrivilegedPlugin_setup_ramWrite_ready) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_TRAP;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        if(PrivilegedPlugin_setup_ramWrite_ready) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        if(PrivilegedPlugin_setup_ramRead_ready) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_XRET;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        if(PrivilegedPlugin_setup_ramRead_ready) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
        PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_IDLE;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
        PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
        PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_IDLE;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_IDLE;
      end
      default : begin
      end
    endcase
    if(PrivilegedPlugin_logic_fsm_wantStart) begin
      PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_IDLE;
    end
    if(PrivilegedPlugin_logic_fsm_wantKill) begin
      PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_BOOT;
    end
  end

  assign when_PrivilegedPlugin_l773 = ((! PrivilegedPlugin_logic_reschedule_payload_fromCommit) && PrivilegedPlugin_logic_decoderInterrupt_raised);
  always @(*) begin
    _zz_PrivilegedPlugin_setup_ramWrite_address = 3'b101;
    case(PrivilegedPlugin_logic_fsm_trap_targetPrivilege)
      2'b01 : begin
        _zz_PrivilegedPlugin_setup_ramWrite_address = 3'b001;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_PrivilegedPlugin_setup_ramWrite_address_1 = 3'b110;
    case(PrivilegedPlugin_logic_fsm_trap_targetPrivilege)
      2'b01 : begin
        _zz_PrivilegedPlugin_setup_ramWrite_address_1 = 3'b010;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_PrivilegedPlugin_setup_ramRead_address = 3'b101;
    case(PrivilegedPlugin_logic_fsm_xret_sourcePrivilege)
      2'b01 : begin
        _zz_PrivilegedPlugin_setup_ramRead_address = 3'b001;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_PrivilegedPlugin_setup_ramRead_address_1 = 3'b111;
    case(PrivilegedPlugin_logic_fsm_trap_targetPrivilege)
      2'b01 : begin
        _zz_PrivilegedPlugin_setup_ramRead_address_1 = 3'b011;
      end
      default : begin
      end
    endcase
  end

  assign when_PrivilegedPlugin_l959 = (PrivilegedPlugin_logic_fsm_xret_targetPrivilege < 2'b11);
  assign switch_PrivilegedPlugin_l960 = PrivilegedPlugin_logic_reschedule_payload_tval[1 : 0];
  assign when_StateMachine_l253_2 = ((! (PrivilegedPlugin_logic_fsm_stateReg == PrivilegedPlugin_logic_fsm_enumDef_IDLE)) && (PrivilegedPlugin_logic_fsm_stateNext == PrivilegedPlugin_logic_fsm_enumDef_IDLE));
  assign CommitPlugin_logic_free_lineEventStream_fifo_io_flush = 1'b0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      HistoryPlugin_logic_update_pushes_2_state <= 24'h000000;
      HistoryPlugin_logic_update_pushes_0_state <= 24'h000000;
      PrivilegedPlugin_setup_privilege <= 2'b11;
      FetchPlugin_stages_1_FETCH_ID <= 12'h000;
      _zz_FetchPlugin_stages_1_isFirstCycle <= 1'b0;
      FetchCachePlugin_logic_invalidate_requested <= 1'b0;
      FetchCachePlugin_logic_invalidate_counter <= 3'b000;
      FetchCachePlugin_logic_invalidate_firstEver <= 1'b1;
      FetchCachePlugin_logic_invalidate_done_regNext <= 1'b0;
      FetchCachePlugin_logic_refill_valid <= 1'b0;
      FetchCachePlugin_logic_refill_hadError <= 1'b0;
      FetchCachePlugin_logic_refill_pushCounter <= 32'h00000000;
      FetchCachePlugin_logic_refill_cmdSent <= 1'b0;
      FetchCachePlugin_logic_refill_wordIndex <= 4'b0000;
      AlignerPlugin_logic_buffer_mask <= 1'b0;
      AlignerPlugin_logic_correctionSent <= 1'b0;
      BranchContextPlugin_logic_ptr_alloc <= 3'b000;
      BranchContextPlugin_logic_ptr_commited <= 3'b000;
      BranchContextPlugin_logic_ptr_free <= 3'b000;
      HistoryPlugin_logic_onCommit_value <= 24'h000000;
      DecoderPredictionPlugin_logic_ras_ptr_push <= 4'b0000;
      DecoderPredictionPlugin_logic_ras_ptr_pop <= 4'b1111;
      BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      _zz_DataCachePlugin_logic_load_ohHistory_1 <= 2'b00;
      _zz_DataCachePlugin_logic_load_ohHistory_2 <= 2'b00;
      CommitPlugin_logic_ptr_alloc <= 5'h00;
      CommitPlugin_logic_ptr_commit <= 5'h00;
      CommitPlugin_logic_ptr_free <= 5'h00;
      CommitPlugin_logic_ptr_empty <= 1'b1;
      CommitPlugin_logic_reschedule_fresh <= 1'b0;
      CommitPlugin_logic_reschedule_valid <= 1'b0;
      CommitPlugin_logic_commit_mask <= 1'b1;
      CommitDebugFilterPlugin_logic_filters_0_value <= 32'h00000000;
      CommitDebugFilterPlugin_logic_filters_1_value <= 32'h00000000;
      CommitDebugFilterPlugin_logic_filters_2_value <= 32'h00000000;
      PrivilegedPlugin_logic_machine_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_machine_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_machine_mstatus_mie <= 1'b0;
      PrivilegedPlugin_logic_machine_mstatus_mpie <= 1'b0;
      PrivilegedPlugin_logic_machine_mstatus_mpp <= 2'b00;
      PrivilegedPlugin_logic_machine_mstatus_fs <= 2'b00;
      PrivilegedPlugin_logic_machine_mstatus_tsr <= 1'b0;
      PrivilegedPlugin_logic_machine_mstatus_tvm <= 1'b0;
      PrivilegedPlugin_logic_machine_mstatus_tw <= 1'b0;
      PrivilegedPlugin_logic_machine_mip_meip <= 1'b0;
      PrivilegedPlugin_logic_machine_mip_mtip <= 1'b0;
      PrivilegedPlugin_logic_machine_mip_msip <= 1'b0;
      PrivilegedPlugin_logic_machine_mie_meie <= 1'b0;
      PrivilegedPlugin_logic_machine_mie_mtie <= 1'b0;
      PrivilegedPlugin_logic_machine_mie_msie <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_iam <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_bp <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_eu <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_es <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_ipf <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_lpf <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_spf <= 1'b0;
      PrivilegedPlugin_logic_machine_mideleg_st <= 1'b0;
      PrivilegedPlugin_logic_machine_mideleg_se <= 1'b0;
      PrivilegedPlugin_logic_machine_mideleg_ss <= 1'b0;
      PrivilegedPlugin_logic_supervisor_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_supervisor_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_supervisor_sstatus_sie <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sstatus_spie <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sstatus_spp <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sip_seipSoft <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sip_stip <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sip_ssip <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sie_seie <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sie_stie <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sie_ssie <= 1'b0;
      PrivilegedPlugin_logic_rescheduleUnbuffered_rValid <= 1'b0;
      EU0_DivPlugin_logic_feed_cmdSent <= 1'b0;
      AguPlugin_logic_fired <= 1'b0;
      LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_0 <= 1'b1;
      LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_0 <= 1'b1;
      DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      DataCachePlugin_mem_toAxi4_awRaw_payload_first <= 1'b1;
      DataCachePlugin_mem_toAxi4_awFiltred_rValid <= 1'b0;
      integer_RfTranslationPlugin_logic_init_counter <= 6'h00;
      integer_RfAllocationPlugin_logic_init_counter <= 7'h01;
      HistoryPlugin_logic_onFetch_value <= 24'h000000;
      Lsu2Plugin_logic_lq_regs_0_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_ptr_priority <= 7'h00;
      Lsu2Plugin_logic_lq_ptr_alloc <= 4'b0000;
      Lsu2Plugin_logic_lq_ptr_free <= 4'b0000;
      Lsu2Plugin_logic_lq_tracker_free <= 4'b1000;
      Lsu2Plugin_logic_lq_reservation_valid <= 1'b0;
      Lsu2Plugin_logic_lq_reservation_counter <= 7'h00;
      Lsu2Plugin_logic_sq_regs_0_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_0_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_0_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_1_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_1_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_1_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_2_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_2_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_2_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_3_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_3_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_3_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_4_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_4_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_4_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_5_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_5_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_5_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_6_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_6_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_6_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_7_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_7_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_7_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_ptr_priority <= 7'h00;
      Lsu2Plugin_logic_sq_ptr_alloc <= 4'b0000;
      Lsu2Plugin_logic_sq_ptr_commit <= 4'b0000;
      Lsu2Plugin_logic_sq_ptr_writeBack <= 4'b0000;
      Lsu2Plugin_logic_sq_ptr_free <= 4'b0000;
      Lsu2Plugin_logic_sq_ptr_onFreeLast_valid <= 1'b0;
      Lsu2Plugin_logic_sq_tracker_free <= 4'b1000;
      Lsu2Plugin_logic_sharedPip_speculativeHitPredictionGotReschedule <= 1'b0;
      Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled <= 1'b1;
      Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask <= 1'b1;
      Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask <= 1'b1;
      Lsu2Plugin_logic_writeback_generation <= 1'b0;
      Lsu2Plugin_logic_writeback_waitOn_refillSlot <= 2'b00;
      Lsu2Plugin_logic_writeback_waitOn_refillSlotAny <= 1'b0;
      toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rValid <= 1'b0;
      Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_valid <= 1'b0;
      Lsu2Plugin_logic_flush_busy <= 1'b0;
      Lsu2Plugin_logic_flush_doit <= 1'b0;
      LsuPlugin_peripheralBus_rsp_valid_regNext <= 1'b0;
      Lsu2Plugin_logic_special_enabled <= 1'b0;
      Lsu2Plugin_logic_special_cmdSent <= 1'b0;
      Lsu2Plugin_logic_special_atomic_lockDelayCounter <= 2'b00;
      Lsu2Plugin_logic_special_atomic_comp_wakeRf <= 1'b0;
      Lsu2Plugin_logic_special_atomic_comp_rfWrite <= 1'b0;
      MmuPlugin_logic_satp_mode <= 1'b0;
      MmuPlugin_logic_satp_ppn <= 20'h00000;
      MmuPlugin_logic_status_mxr <= 1'b0;
      MmuPlugin_logic_status_sum <= 1'b0;
      MmuPlugin_logic_status_mprv <= 1'b0;
      FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value <= 2'b00;
      FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value <= 1'b0;
      Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value <= 2'b00;
      Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value <= 1'b0;
      Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg <= 1'b1;
      Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg <= 1'b1;
      CsrRamPlugin_logic_flush_counter <= 4'b0000;
      PrivilegedPlugin_logic_decoderInterrupt_raised <= 1'b0;
      PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt <= 1'b0;
      PrivilegedPlugin_logic_decoderInterrupt_counter <= 3'b000;
      EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired <= 1'b0;
      EU0_CsrAccessPlugin_logic_fsm_stateReg <= EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT;
      EnvCallPlugin_logic_flushes_stateReg <= EnvCallPlugin_logic_flushes_enumDef_BOOT;
      FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg <= 1'b1;
      MmuPlugin_logic_refill_cacheRefill <= 2'b00;
      MmuPlugin_logic_refill_cacheRefillAny <= 1'b0;
      MmuPlugin_logic_refill_load_rsp_valid <= 1'b0;
      MmuPlugin_logic_invalidate_requested <= 1'b1;
      MmuPlugin_logic_invalidate_counter <= 3'b000;
      MmuPlugin_logic_invalidate_done_regNext <= 1'b0;
      Lsu2Plugin_logic_sharedPip_stages_1_valid <= 1'b0;
      Lsu2Plugin_logic_sharedPip_stages_2_valid <= 1'b0;
      Lsu2Plugin_logic_sharedPip_stages_3_valid <= 1'b0;
      Lsu2Plugin_logic_lqSqArbitration_s1_valid <= 1'b0;
      Lsu2Plugin_logic_special_atomic_stateReg <= Lsu2Plugin_logic_special_atomic_enumDef_BOOT;
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_enumDef_BOOT;
      DecoderPlugin_logic_exception_trigged <= 1'b0;
      DecoderPlugin_logic_exception_doItAgain <= 1'b0;
      FrontendPlugin_decoded_OP_ID <= 12'h000;
      DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle <= 1'b1;
      ALU0_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      EU0_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      EU0_ExecutionUnitBase_pipeline_execute_1_valid <= 1'b0;
      EU0_ExecutionUnitBase_pipeline_execute_2_valid <= 1'b0;
      DispatchPlugin_logic_ptr_next <= 4'b1001;
      DispatchPlugin_logic_ptr_current <= 4'b1000;
      DispatchPlugin_logic_push_fenceYoungerLast <= 1'b0;
      DispatchPlugin_logic_pop_0_stagesList_1_valid <= 1'b0;
      DispatchPlugin_logic_pop_1_stagesList_1_valid <= 1'b0;
      RfDependencyPlugin_logic_forRf_integer_init_counter <= 7'h00;
      FrontendPlugin_dispatch_valid <= 1'b0;
      FrontendPlugin_serialized_valid <= 1'b0;
      PcPlugin_logic_init_counter <= 7'h00;
      PcPlugin_logic_fetchPc_pcReg <= externalResetVector;
      PcPlugin_logic_fetchPc_correctionReg <= 1'b0;
      PcPlugin_logic_fetchPc_inc <= 1'b0;
      FetchPlugin_stages_1_valid <= 1'b0;
      FetchPlugin_stages_2_valid <= 1'b0;
      FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid <= 1'b0;
      PrivilegedPlugin_logic_fsm_stateReg <= PrivilegedPlugin_logic_fsm_enumDef_BOOT;
    end else begin
      FetchPlugin_stages_1_FETCH_ID <= (FetchPlugin_stages_1_FETCH_ID + _zz_FetchPlugin_stages_1_FETCH_ID);
      if(FetchPlugin_stages_1_valid) begin
        _zz_FetchPlugin_stages_1_isFirstCycle <= 1'b1;
      end
      if(when_Stage_l170) begin
        _zz_FetchPlugin_stages_1_isFirstCycle <= 1'b0;
      end
      if(FetchCachePlugin_setup_invalidatePort_cmd_valid) begin
        FetchCachePlugin_logic_invalidate_requested <= 1'b1;
      end
      if(FetchCachePlugin_logic_invalidate_done) begin
        FetchCachePlugin_logic_invalidate_firstEver <= 1'b0;
      end
      if(when_FetchCachePlugin_l379) begin
        FetchCachePlugin_logic_invalidate_counter <= (FetchCachePlugin_logic_invalidate_counter + 3'b001);
      end
      if(when_FetchCachePlugin_l391) begin
        FetchCachePlugin_logic_invalidate_counter <= 3'b000;
        FetchCachePlugin_logic_invalidate_requested <= 1'b0;
      end
      FetchCachePlugin_logic_invalidate_done_regNext <= FetchCachePlugin_logic_invalidate_done;
      if(FetchCachePlugin_logic_refill_fire) begin
        FetchCachePlugin_logic_refill_valid <= 1'b0;
      end
      if(when_FetchCachePlugin_l422) begin
        if(FetchCachePlugin_logic_refill_start_valid) begin
          FetchCachePlugin_logic_refill_valid <= 1'b1;
          FetchCachePlugin_logic_refill_pushCounter <= (FetchCachePlugin_logic_refill_pushCounter + 32'h00000001);
        end
      end
      if(FetchCachePlugin_mem_cmd_fire) begin
        FetchCachePlugin_logic_refill_cmdSent <= 1'b1;
      end
      if(FetchCachePlugin_logic_refill_fire) begin
        FetchCachePlugin_logic_refill_cmdSent <= 1'b0;
      end
      if(FetchCachePlugin_mem_rsp_valid) begin
        FetchCachePlugin_logic_refill_wordIndex <= (FetchCachePlugin_logic_refill_wordIndex + 4'b0001);
        if(FetchCachePlugin_mem_rsp_payload_error) begin
          FetchCachePlugin_logic_refill_hadError <= 1'b1;
        end
      end
      if(FetchCachePlugin_logic_refill_fire) begin
        FetchCachePlugin_logic_refill_hadError <= 1'b0;
      end
      if(AlignerPlugin_logic_fireOutput) begin
        AlignerPlugin_logic_buffer_mask <= AlignerPlugin_logic_slices_remains_1[0 : 0];
      end
      if(AlignerPlugin_logic_fireInput) begin
        AlignerPlugin_logic_buffer_mask <= ((AlignerPlugin_logic_fireOutput ? AlignerPlugin_logic_slices_remains_1[1 : 1] : AlignerPlugin_setup_s2m_MASK_FRONT) & AlignerPlugin_logic_postMask);
      end
      if(AlignerPlugin_setup_sequenceJump_valid) begin
        AlignerPlugin_logic_correctionSent <= 1'b1;
      end
      if(when_AlignerPlugin_l264) begin
        AlignerPlugin_logic_correctionSent <= 1'b0;
      end
      if(FrontendPlugin_aligned_isFlushed) begin
        AlignerPlugin_logic_buffer_mask <= 1'b0;
      end
      if(FrontendPlugin_allocated_isFireing) begin
        BranchContextPlugin_logic_ptr_alloc <= BranchContextPlugin_logic_alloc_allocNext_1;
      end
      DecoderPredictionPlugin_logic_ras_ptr_push <= (_zz_DecoderPredictionPlugin_logic_ras_ptr_push - _zz_DecoderPredictionPlugin_logic_ras_ptr_push_3);
      DecoderPredictionPlugin_logic_ras_ptr_pop <= (_zz_DecoderPredictionPlugin_logic_ras_ptr_pop - _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_3);
      if(FetchPlugin_stages_1_valid) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b1;
      end
      if(when_BtbPlugin_l109) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      end
      _zz_DataCachePlugin_logic_load_ohHistory_1 <= _zz_DataCachePlugin_logic_load_ohHistory_0;
      _zz_DataCachePlugin_logic_load_ohHistory_2 <= _zz_DataCachePlugin_logic_load_ohHistory_1;
      CommitPlugin_logic_ptr_commit <= CommitPlugin_logic_ptr_commitNext;
      CommitPlugin_logic_ptr_alloc <= CommitPlugin_logic_ptr_allocNext;
      CommitPlugin_logic_ptr_empty <= (CommitPlugin_logic_ptr_allocNext == CommitPlugin_logic_ptr_commitNext);
      CommitPlugin_logic_reschedule_fresh <= 1'b0;
      if(when_CommitPlugin_l131) begin
        CommitPlugin_logic_reschedule_fresh <= 1'b1;
        CommitPlugin_logic_reschedule_valid <= 1'b1;
      end
      CommitPlugin_logic_commit_mask <= CommitPlugin_logic_commit_maskComb;
      if(CommitPlugin_logic_commit_rescheduleHit) begin
        CommitPlugin_logic_reschedule_valid <= 1'b0;
      end
      if(when_CommitPlugin_l194) begin
        if(when_CommitPlugin_l217) begin
          CommitPlugin_logic_commit_mask <= 1'b1;
        end
      end
      if(CommitPlugin_logic_ptr_canFree) begin
        CommitPlugin_logic_ptr_free <= (CommitPlugin_logic_ptr_free + 5'h01);
      end
      CommitDebugFilterPlugin_logic_filters_0_value <= (CommitDebugFilterPlugin_logic_filters_0_value + _zz_CommitDebugFilterPlugin_logic_filters_0_value);
      CommitDebugFilterPlugin_logic_filters_1_value <= (CommitDebugFilterPlugin_logic_filters_1_value + _zz_CommitDebugFilterPlugin_logic_filters_1_value);
      CommitDebugFilterPlugin_logic_filters_2_value <= (CommitDebugFilterPlugin_logic_filters_2_value + _zz_CommitDebugFilterPlugin_logic_filters_2_value);
      PrivilegedPlugin_logic_machine_mip_meip <= PrivilegedPlugin_io_int_machine_external;
      PrivilegedPlugin_logic_machine_mip_mtip <= PrivilegedPlugin_io_int_machine_timer;
      PrivilegedPlugin_logic_machine_mip_msip <= PrivilegedPlugin_io_int_machine_software;
      if(PrivilegedPlugin_logic_rescheduleUnbuffered_ready) begin
        PrivilegedPlugin_logic_rescheduleUnbuffered_rValid <= PrivilegedPlugin_logic_rescheduleUnbuffered_valid;
      end
      if(toplevel_EU0_DivPlugin_logic_div_io_cmd_fire) begin
        EU0_DivPlugin_logic_feed_cmdSent <= 1'b1;
      end
      if(when_DivPlugin_l76) begin
        EU0_DivPlugin_logic_feed_cmdSent <= 1'b0;
      end
      if(AguPlugin_setup_port_valid) begin
        AguPlugin_logic_fired <= 1'b1;
      end
      if(when_AguPlugin_l89) begin
        AguPlugin_logic_fired <= 1'b0;
      end
      if(LsuPlugin_peripheralBus_toAxiLite4_a_fire) begin
        LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(LsuPlugin_peripheralBus_toAxiLite4_wRaw_fire) begin
        LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(LsuPlugin_peripheralBus_cmd_ready) begin
        LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_0 <= 1'b1;
        LsuPlugin_peripheralBus_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(DataCachePlugin_mem_toAxi4_awRaw_fire) begin
        DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(DataCachePlugin_mem_toAxi4_wRaw_fire) begin
        DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(DataCachePlugin_mem_write_cmd_ready) begin
        DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_0 <= 1'b1;
        DataCachePlugin_mem_write_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(DataCachePlugin_mem_toAxi4_awRaw_fire) begin
        DataCachePlugin_mem_toAxi4_awRaw_payload_first <= DataCachePlugin_mem_toAxi4_awRaw_payload_last;
      end
      if(DataCachePlugin_mem_toAxi4_awFiltred_ready) begin
        DataCachePlugin_mem_toAxi4_awFiltred_rValid <= DataCachePlugin_mem_toAxi4_awFiltred_valid;
      end
      if(integer_RfTranslationPlugin_logic_init_busy) begin
        integer_RfTranslationPlugin_logic_init_counter <= (integer_RfTranslationPlugin_logic_init_counter + 6'h01);
      end
      if(integer_RfAllocationPlugin_logic_init_busy) begin
        integer_RfAllocationPlugin_logic_init_counter <= (integer_RfAllocationPlugin_logic_init_counter + 7'h01);
      end
      BranchContextPlugin_logic_ptr_commited <= BranchContextPlugin_logic_onCommit_commitedNext;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        BranchContextPlugin_logic_ptr_alloc <= BranchContextPlugin_logic_onCommit_commitedNext;
      end
      HistoryPlugin_logic_onCommit_value <= HistoryPlugin_logic_onCommit_valueNext_1;
      HistoryPlugin_logic_onFetch_value <= HistoryPlugin_logic_onFetch_valueNext;
      HistoryPlugin_logic_update_pushes_0_state <= HistoryPlugin_logic_update_pushes_0_stateNext_1;
      if(FetchCachePlugin_setup_historyJump_valid) begin
        HistoryPlugin_logic_update_pushes_0_state <= FetchCachePlugin_setup_historyJump_payload_history;
      end
      HistoryPlugin_logic_update_pushes_2_state <= HistoryPlugin_logic_update_pushes_2_stateNext_1;
      if(DecoderPredictionPlugin_setup_historyPush_flush) begin
        HistoryPlugin_logic_update_pushes_0_state <= HistoryPlugin_logic_update_pushes_2_stateNext_1;
      end
      if(CommitPlugin_logic_reschedule_reschedulePort_valid) begin
        HistoryPlugin_logic_update_pushes_2_state <= HistoryPlugin_logic_update_rescheduleFlush_newHistory;
        HistoryPlugin_logic_update_pushes_0_state <= HistoryPlugin_logic_update_rescheduleFlush_newHistory;
      end
      if(CommitPlugin_logic_reschedule_reschedulePort_valid) begin
        DecoderPredictionPlugin_logic_ras_ptr_push <= DecoderPredictionPlugin_logic_ras_healPush;
        DecoderPredictionPlugin_logic_ras_ptr_pop <= DecoderPredictionPlugin_logic_ras_healPop;
      end
      Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_0_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_0_allocation) begin
        Lsu2Plugin_logic_lq_regs_0_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_0_redoSet) begin
        Lsu2Plugin_logic_lq_regs_0_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_0_delete) begin
        Lsu2Plugin_logic_lq_regs_0_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_0_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338) begin
        Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_1_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_1_allocation) begin
        Lsu2Plugin_logic_lq_regs_1_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_1_redoSet) begin
        Lsu2Plugin_logic_lq_regs_1_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_1_delete) begin
        Lsu2Plugin_logic_lq_regs_1_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_1_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_1) begin
        Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_2_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_2_allocation) begin
        Lsu2Plugin_logic_lq_regs_2_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_2_redoSet) begin
        Lsu2Plugin_logic_lq_regs_2_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_2_delete) begin
        Lsu2Plugin_logic_lq_regs_2_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_2_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_2) begin
        Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_3_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_3_allocation) begin
        Lsu2Plugin_logic_lq_regs_3_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_3_redoSet) begin
        Lsu2Plugin_logic_lq_regs_3_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_3_delete) begin
        Lsu2Plugin_logic_lq_regs_3_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_3_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_3) begin
        Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_4_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_4_allocation) begin
        Lsu2Plugin_logic_lq_regs_4_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_4_redoSet) begin
        Lsu2Plugin_logic_lq_regs_4_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_4_delete) begin
        Lsu2Plugin_logic_lq_regs_4_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_4_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_4) begin
        Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_5_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_5_allocation) begin
        Lsu2Plugin_logic_lq_regs_5_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_5_redoSet) begin
        Lsu2Plugin_logic_lq_regs_5_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_5_delete) begin
        Lsu2Plugin_logic_lq_regs_5_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_5_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_5) begin
        Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_6_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_6_allocation) begin
        Lsu2Plugin_logic_lq_regs_6_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_6_redoSet) begin
        Lsu2Plugin_logic_lq_regs_6_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_6_delete) begin
        Lsu2Plugin_logic_lq_regs_6_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_6_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_6) begin
        Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_7_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_7_allocation) begin
        Lsu2Plugin_logic_lq_regs_7_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_7_redoSet) begin
        Lsu2Plugin_logic_lq_regs_7_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_7_delete) begin
        Lsu2Plugin_logic_lq_regs_7_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_7_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_7) begin
        Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_tracker_free <= Lsu2Plugin_logic_lq_tracker_freeNext;
      Lsu2Plugin_logic_lq_ptr_priority <= Lsu2Plugin_logic_lq_onCommit_priority_1;
      Lsu2Plugin_logic_lq_ptr_free <= (Lsu2Plugin_logic_lq_ptr_free + _zz_Lsu2Plugin_logic_lq_ptr_free);
      if(Lsu2Plugin_logic_lq_reservation_kill) begin
        Lsu2Plugin_logic_lq_reservation_valid <= 1'b0;
      end
      if(when_Lsu2Plugin_l484) begin
        Lsu2Plugin_logic_lq_reservation_valid <= 1'b0;
      end else begin
        Lsu2Plugin_logic_lq_reservation_counter <= (Lsu2Plugin_logic_lq_reservation_counter + 7'h01);
      end
      Lsu2Plugin_logic_sq_regs_0_commited <= Lsu2Plugin_logic_sq_regs_0_commitedNext;
      Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_0_allocation) begin
        Lsu2Plugin_logic_sq_regs_0_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_0_redoSet) begin
        Lsu2Plugin_logic_sq_regs_0_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_0_delete) begin
        Lsu2Plugin_logic_sq_regs_0_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_0_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_0_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385) begin
        Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_1_commited <= Lsu2Plugin_logic_sq_regs_1_commitedNext;
      Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_1_allocation) begin
        Lsu2Plugin_logic_sq_regs_1_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_1_redoSet) begin
        Lsu2Plugin_logic_sq_regs_1_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_1_delete) begin
        Lsu2Plugin_logic_sq_regs_1_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_1_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_1_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_1) begin
        Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_2_commited <= Lsu2Plugin_logic_sq_regs_2_commitedNext;
      Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_2_allocation) begin
        Lsu2Plugin_logic_sq_regs_2_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_2_redoSet) begin
        Lsu2Plugin_logic_sq_regs_2_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_2_delete) begin
        Lsu2Plugin_logic_sq_regs_2_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_2_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_2_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_2) begin
        Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_3_commited <= Lsu2Plugin_logic_sq_regs_3_commitedNext;
      Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_3_allocation) begin
        Lsu2Plugin_logic_sq_regs_3_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_3_redoSet) begin
        Lsu2Plugin_logic_sq_regs_3_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_3_delete) begin
        Lsu2Plugin_logic_sq_regs_3_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_3_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_3_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_3) begin
        Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_4_commited <= Lsu2Plugin_logic_sq_regs_4_commitedNext;
      Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_4_allocation) begin
        Lsu2Plugin_logic_sq_regs_4_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_4_redoSet) begin
        Lsu2Plugin_logic_sq_regs_4_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_4_delete) begin
        Lsu2Plugin_logic_sq_regs_4_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_4_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_4_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_4) begin
        Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_5_commited <= Lsu2Plugin_logic_sq_regs_5_commitedNext;
      Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_5_allocation) begin
        Lsu2Plugin_logic_sq_regs_5_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_5_redoSet) begin
        Lsu2Plugin_logic_sq_regs_5_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_5_delete) begin
        Lsu2Plugin_logic_sq_regs_5_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_5_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_5_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_5) begin
        Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_6_commited <= Lsu2Plugin_logic_sq_regs_6_commitedNext;
      Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_6_allocation) begin
        Lsu2Plugin_logic_sq_regs_6_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_6_redoSet) begin
        Lsu2Plugin_logic_sq_regs_6_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_6_delete) begin
        Lsu2Plugin_logic_sq_regs_6_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_6_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_6_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_6) begin
        Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_7_commited <= Lsu2Plugin_logic_sq_regs_7_commitedNext;
      Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_7_allocation) begin
        Lsu2Plugin_logic_sq_regs_7_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_7_redoSet) begin
        Lsu2Plugin_logic_sq_regs_7_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_7_delete) begin
        Lsu2Plugin_logic_sq_regs_7_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_7_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_7_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_7) begin
        Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_ptr_commit <= Lsu2Plugin_logic_sq_ptr_commitNext;
      Lsu2Plugin_logic_sq_ptr_onFreeLast_valid <= Lsu2Plugin_logic_sq_ptr_onFree_valid;
      Lsu2Plugin_logic_sq_tracker_free <= Lsu2Plugin_logic_sq_tracker_freeNext;
      if(FrontendPlugin_dispatch_isFireing) begin
        Lsu2Plugin_logic_lq_ptr_alloc <= Lsu2Plugin_logic_allocation_loads_alloc_1;
        Lsu2Plugin_logic_sq_ptr_alloc <= Lsu2Plugin_logic_allocation_stores_alloc_1;
      end
      if(Lsu2Plugin_logic_lqSqArbitration_s0_ready) begin
        if(Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT) begin
          if(Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[0]) begin
            Lsu2Plugin_logic_lq_regs_0_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID) begin
            Lsu2Plugin_logic_lq_regs_1_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_1) begin
            Lsu2Plugin_logic_lq_regs_2_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2) begin
            Lsu2Plugin_logic_lq_regs_3_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_3) begin
            Lsu2Plugin_logic_lq_regs_4_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4) begin
            Lsu2Plugin_logic_lq_regs_5_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5) begin
            Lsu2Plugin_logic_lq_regs_6_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6) begin
            Lsu2Plugin_logic_lq_regs_7_redo <= 1'b0;
          end
        end
        if(Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT) begin
          if(Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[0]) begin
            Lsu2Plugin_logic_sq_regs_0_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID) begin
            Lsu2Plugin_logic_sq_regs_1_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_1) begin
            Lsu2Plugin_logic_sq_regs_2_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2) begin
            Lsu2Plugin_logic_sq_regs_3_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_3) begin
            Lsu2Plugin_logic_sq_regs_4_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4) begin
            Lsu2Plugin_logic_sq_regs_5_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5) begin
            Lsu2Plugin_logic_sq_regs_6_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6) begin
            Lsu2Plugin_logic_sq_regs_7_redo <= 1'b0;
          end
        end
      end
      if(Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap) begin
        Lsu2Plugin_logic_sharedPip_speculativeHitPredictionGotReschedule <= 1'b0;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_sharedPip_speculativeHitPredictionGotReschedule <= 1'b1;
      end
      if(Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap) begin
        Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled <= 1'b0;
      end
      if(Lsu2Plugin_logic_sharedPip_speculateHitTrapRecovered) begin
        Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled <= 1'b1;
      end
      if(when_Lsu2Plugin_l841) begin
        if(when_Lsu2Plugin_l843) begin
          if(Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ) begin
            Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask <= 1'b0;
          end
          if(when_Lsu2Plugin_l845) begin
            Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask <= 1'b0;
          end
        end
      end
      if(when_Lsu2Plugin_l849) begin
        Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask <= 1'b1;
        Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask <= 1'b1;
      end
      if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
        case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
          Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
          end
          Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          end
          Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
          end
          Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          end
          Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          end
          Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
          end
          Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
          end
          default : begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
              if(when_Lsu2Plugin_l1333) begin
                if(Lsu2Plugin_logic_sharedPip_stages_3_LR) begin
                  Lsu2Plugin_logic_lq_reservation_valid <= (! Lsu2Plugin_logic_lq_reservation_valid);
                  Lsu2Plugin_logic_lq_reservation_counter <= 7'h00;
                end
              end
            end
          end
        endcase
      end
      Lsu2Plugin_logic_writeback_waitOn_refillSlot <= ((Lsu2Plugin_logic_writeback_waitOn_refillSlot | Lsu2Plugin_logic_writeback_waitOn_refillSlotSet) & (~ DataCachePlugin_setup_refillCompletions));
      Lsu2Plugin_logic_writeback_waitOn_refillSlotAny <= ((Lsu2Plugin_logic_writeback_waitOn_refillSlotAny || Lsu2Plugin_logic_writeback_waitOn_refillSlotAnySet) && (! (|DataCachePlugin_setup_refillCompletions)));
      if(Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready) begin
        toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rValid <= Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_valid;
      end
      Lsu2Plugin_logic_sq_ptr_writeBack <= (Lsu2Plugin_logic_sq_ptr_writeBack + _zz_Lsu2Plugin_logic_sq_ptr_writeBack);
      Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_valid <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_valid;
      if(when_Lsu2Plugin_l1488) begin
        if(Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
          Lsu2Plugin_logic_writeback_generation <= (! Lsu2Plugin_logic_writeback_generation);
          Lsu2Plugin_logic_sq_ptr_writeBack <= Lsu2Plugin_logic_sq_ptr_free;
        end
      end
      if(when_Lsu2Plugin_l1509) begin
        Lsu2Plugin_logic_sq_ptr_writeBack <= (Lsu2Plugin_logic_sq_ptr_writeBack + 4'b0001);
      end
      if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
        Lsu2Plugin_logic_sq_ptr_free <= (Lsu2Plugin_logic_sq_ptr_free + 4'b0001);
        Lsu2Plugin_logic_sq_ptr_priority <= (Lsu2Plugin_logic_sq_ptr_priority <<< 1);
        if(when_Lsu2Plugin_l1521) begin
          Lsu2Plugin_logic_sq_ptr_priority <= 7'h7f;
        end
      end
      Lsu2Plugin_logic_flush_doit <= (Lsu2Plugin_logic_sq_ptr_commit == Lsu2Plugin_logic_sq_ptr_free);
      if(Lsu2Plugin_setup_flushPort_cmd_valid) begin
        Lsu2Plugin_logic_flush_busy <= 1'b1;
        Lsu2Plugin_logic_flush_doit <= 1'b0;
      end
      if(when_Lsu2Plugin_l1553) begin
        if(when_Lsu2Plugin_l1561) begin
          if(Lsu2Plugin_setup_cacheStore_rsp_payload_redo) begin
            Lsu2Plugin_logic_writeback_generation <= (! Lsu2Plugin_logic_writeback_generation);
          end
        end
        if(when_Lsu2Plugin_l1569) begin
          Lsu2Plugin_logic_flush_busy <= 1'b0;
        end
      end
      LsuPlugin_peripheralBus_rsp_valid_regNext <= LsuPlugin_peripheralBus_rsp_valid;
      if(Lsu2Plugin_logic_special_hit) begin
        Lsu2Plugin_logic_special_enabled <= 1'b1;
      end
      if(Lsu2Plugin_logic_special_fire) begin
        Lsu2Plugin_logic_special_enabled <= 1'b0;
      end
      if(LsuPlugin_peripheralBus_cmd_fire) begin
        Lsu2Plugin_logic_special_cmdSent <= 1'b1;
      end
      if(Lsu2Plugin_logic_special_fire) begin
        Lsu2Plugin_logic_special_cmdSent <= 1'b0;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_lq_ptr_free <= 4'b0000;
        Lsu2Plugin_logic_lq_ptr_alloc <= 4'b0000;
        Lsu2Plugin_logic_lq_ptr_priority <= 7'h00;
        Lsu2Plugin_logic_sq_ptr_alloc <= Lsu2Plugin_logic_sq_ptr_commitNext;
        Lsu2Plugin_logic_special_enabled <= 1'b0;
      end
      if(PrivilegedPlugin_setup_xretAwayFromMachine) begin
        MmuPlugin_logic_status_mprv <= 1'b0;
      end
      FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value <= FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
      FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value <= FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_valueNext;
      Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value <= Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
      Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value <= Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_valueNext;
      Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg <= Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL_overloaded;
      if(when_MmuPlugin_l278) begin
        Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg <= 1'b1;
      end
      Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg <= Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded;
      if(when_MmuPlugin_l278_1) begin
        Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg <= 1'b1;
      end
      if(when_CsrRamPlugin_l61) begin
        CsrRamPlugin_logic_flush_counter <= (CsrRamPlugin_logic_flush_counter + 4'b0001);
      end
      PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt <= PrivilegedPlugin_logic_interrupt_valid;
      if(PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt) begin
        PrivilegedPlugin_logic_decoderInterrupt_counter <= (PrivilegedPlugin_logic_decoderInterrupt_counter + 3'b001);
      end
      if(when_PrivilegedPlugin_l675) begin
        PrivilegedPlugin_logic_decoderInterrupt_counter <= 3'b000;
      end
      if(when_PrivilegedPlugin_l679) begin
        PrivilegedPlugin_logic_decoderInterrupt_raised <= 1'b1;
      end
      if(when_CsrAccessPlugin_l328) begin
        PrivilegedPlugin_logic_machine_cause_interrupt <= EU0_CsrAccessPlugin_setup_onWriteBits[31];
        PrivilegedPlugin_logic_machine_cause_code <= EU0_CsrAccessPlugin_setup_onWriteBits[3 : 0];
      end
      if(when_CsrAccessPlugin_l328_1) begin
        PrivilegedPlugin_logic_machine_mstatus_mpp <= EU0_CsrAccessPlugin_setup_onWriteBits[12 : 11];
        PrivilegedPlugin_logic_machine_mstatus_mpie <= EU0_CsrAccessPlugin_setup_onWriteBits[7];
        PrivilegedPlugin_logic_machine_mstatus_mie <= EU0_CsrAccessPlugin_setup_onWriteBits[3];
        PrivilegedPlugin_logic_machine_mstatus_tsr <= EU0_CsrAccessPlugin_setup_onWriteBits[22];
        PrivilegedPlugin_logic_machine_mstatus_tw <= EU0_CsrAccessPlugin_setup_onWriteBits[21];
        PrivilegedPlugin_logic_machine_mstatus_tvm <= EU0_CsrAccessPlugin_setup_onWriteBits[20];
        PrivilegedPlugin_logic_machine_mstatus_fs <= EU0_CsrAccessPlugin_setup_onWriteBits[14 : 13];
        PrivilegedPlugin_logic_supervisor_sstatus_spp <= EU0_CsrAccessPlugin_setup_onWriteBits[8 : 8];
        PrivilegedPlugin_logic_supervisor_sstatus_spie <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_supervisor_sstatus_sie <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
        MmuPlugin_logic_status_mxr <= EU0_CsrAccessPlugin_setup_onWriteBits[19];
        MmuPlugin_logic_status_sum <= EU0_CsrAccessPlugin_setup_onWriteBits[18];
        MmuPlugin_logic_status_mprv <= EU0_CsrAccessPlugin_setup_onWriteBits[17];
      end
      if(when_CsrAccessPlugin_l328_2) begin
        PrivilegedPlugin_logic_supervisor_sip_seipSoft <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        PrivilegedPlugin_logic_supervisor_sip_stip <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_supervisor_sip_ssip <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
      end
      if(when_CsrAccessPlugin_l328_3) begin
        PrivilegedPlugin_logic_machine_mie_meie <= EU0_CsrAccessPlugin_setup_onWriteBits[11];
        PrivilegedPlugin_logic_machine_mie_mtie <= EU0_CsrAccessPlugin_setup_onWriteBits[7];
        PrivilegedPlugin_logic_machine_mie_msie <= EU0_CsrAccessPlugin_setup_onWriteBits[3];
        PrivilegedPlugin_logic_supervisor_sie_seie <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        PrivilegedPlugin_logic_supervisor_sie_stie <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_supervisor_sie_ssie <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
      end
      if(when_CsrAccessPlugin_l328_4) begin
        PrivilegedPlugin_logic_machine_medeleg_iam <= EU0_CsrAccessPlugin_setup_onWriteBits[0];
        PrivilegedPlugin_logic_machine_medeleg_bp <= EU0_CsrAccessPlugin_setup_onWriteBits[3];
        PrivilegedPlugin_logic_machine_medeleg_eu <= EU0_CsrAccessPlugin_setup_onWriteBits[8];
        PrivilegedPlugin_logic_machine_medeleg_es <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        PrivilegedPlugin_logic_machine_medeleg_ipf <= EU0_CsrAccessPlugin_setup_onWriteBits[12];
        PrivilegedPlugin_logic_machine_medeleg_lpf <= EU0_CsrAccessPlugin_setup_onWriteBits[13];
        PrivilegedPlugin_logic_machine_medeleg_spf <= EU0_CsrAccessPlugin_setup_onWriteBits[15];
      end
      if(when_CsrAccessPlugin_l328_5) begin
        PrivilegedPlugin_logic_machine_mideleg_se <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        PrivilegedPlugin_logic_machine_mideleg_st <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_machine_mideleg_ss <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
      end
      if(when_CsrAccessPlugin_l328_6) begin
        PrivilegedPlugin_logic_supervisor_cause_interrupt <= EU0_CsrAccessPlugin_setup_onWriteBits[31];
        PrivilegedPlugin_logic_supervisor_cause_code <= EU0_CsrAccessPlugin_setup_onWriteBits[3 : 0];
      end
      if(when_CsrAccessPlugin_l328_7) begin
        PrivilegedPlugin_logic_supervisor_sstatus_spp <= EU0_CsrAccessPlugin_setup_onWriteBits[8 : 8];
        PrivilegedPlugin_logic_supervisor_sstatus_spie <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_supervisor_sstatus_sie <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
        PrivilegedPlugin_logic_machine_mstatus_fs <= EU0_CsrAccessPlugin_setup_onWriteBits[14 : 13];
        MmuPlugin_logic_status_mxr <= EU0_CsrAccessPlugin_setup_onWriteBits[19];
        MmuPlugin_logic_status_sum <= EU0_CsrAccessPlugin_setup_onWriteBits[18];
      end
      if(when_CsrAccessPlugin_l328_8) begin
        if(PrivilegedPlugin_logic_machine_mideleg_se) begin
          PrivilegedPlugin_logic_supervisor_sie_seie <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        end
        if(PrivilegedPlugin_logic_machine_mideleg_st) begin
          PrivilegedPlugin_logic_supervisor_sie_stie <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        end
        if(PrivilegedPlugin_logic_machine_mideleg_ss) begin
          PrivilegedPlugin_logic_supervisor_sie_ssie <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
        end
      end
      if(when_CsrAccessPlugin_l328_9) begin
        if(PrivilegedPlugin_logic_machine_mideleg_ss) begin
          PrivilegedPlugin_logic_supervisor_sip_ssip <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
        end
      end
      if(when_CsrAccessPlugin_l333) begin
        if(when_CsrAccessPlugin_l328_10) begin
          MmuPlugin_logic_satp_mode <= EU0_CsrAccessPlugin_setup_onWriteBits[31 : 31];
          MmuPlugin_logic_satp_ppn <= EU0_CsrAccessPlugin_setup_onWriteBits[19 : 0];
        end
      end
      if(when_CsrAccessPlugin_l338) begin
        EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired <= 1'b1;
      end
      if(EU0_CsrAccessPlugin_setup_onWriteMovingOff) begin
        EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired <= 1'b0;
      end
      EU0_CsrAccessPlugin_logic_fsm_stateReg <= EU0_CsrAccessPlugin_logic_fsm_stateNext;
      EnvCallPlugin_logic_flushes_stateReg <= EnvCallPlugin_logic_flushes_stateNext;
      FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg <= FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded;
      if(when_MmuPlugin_l278_2) begin
        FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg <= 1'b1;
      end
      MmuPlugin_logic_refill_cacheRefill <= ((MmuPlugin_logic_refill_cacheRefill | MmuPlugin_logic_refill_cacheRefillSet) & (~ DataCachePlugin_setup_refillCompletions));
      MmuPlugin_logic_refill_cacheRefillAny <= ((MmuPlugin_logic_refill_cacheRefillAny || MmuPlugin_logic_refill_cacheRefillAnySet) && (! (|DataCachePlugin_setup_refillCompletions)));
      MmuPlugin_logic_refill_load_rsp_valid <= MmuPlugin_setup_cacheLoad_rsp_valid;
      if(MmuPlugin_setup_invalidatePort_cmd_valid) begin
        MmuPlugin_logic_invalidate_requested <= 1'b1;
      end
      if(when_MmuPlugin_l522) begin
        MmuPlugin_logic_invalidate_counter <= (MmuPlugin_logic_invalidate_counter + 3'b001);
      end
      if(when_MmuPlugin_l535) begin
        MmuPlugin_logic_invalidate_counter <= 3'b000;
        MmuPlugin_logic_invalidate_requested <= 1'b0;
      end
      MmuPlugin_logic_invalidate_done_regNext <= MmuPlugin_logic_invalidate_done;
      Lsu2Plugin_logic_sharedPip_stages_1_valid <= _zz_Lsu2Plugin_logic_sharedPip_stages_1_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_sharedPip_stages_1_valid <= 1'b0;
      end
      Lsu2Plugin_logic_sharedPip_stages_2_valid <= Lsu2Plugin_logic_sharedPip_stages_1_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_sharedPip_stages_2_valid <= 1'b0;
      end
      Lsu2Plugin_logic_sharedPip_stages_3_valid <= Lsu2Plugin_logic_sharedPip_stages_2_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_sharedPip_stages_3_valid <= 1'b0;
      end
      if(Lsu2Plugin_logic_lqSqArbitration_s0_ready_output) begin
        Lsu2Plugin_logic_lqSqArbitration_s1_valid <= Lsu2Plugin_logic_lqSqArbitration_s0_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_lqSqArbitration_s1_valid <= 1'b0;
      end
      Lsu2Plugin_logic_special_atomic_stateReg <= Lsu2Plugin_logic_special_atomic_stateNext;
      (* parallel_case *)
      case(1) // synthesis parallel_case
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
        end
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
        end
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
          if(Lsu2Plugin_setup_cacheLoad_rsp_valid) begin
            Lsu2Plugin_logic_special_atomic_comp_rfWrite <= 1'b0;
          end
        end
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
          Lsu2Plugin_logic_special_atomic_lockDelayCounter <= (Lsu2Plugin_logic_special_atomic_lockDelayCounter + 2'b01);
        end
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
        end
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
          Lsu2Plugin_logic_special_atomic_comp_wakeRf <= 1'b0;
          Lsu2Plugin_logic_special_atomic_comp_rfWrite <= 1'b0;
        end
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
        end
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
        end
        (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l253) begin
        Lsu2Plugin_logic_special_atomic_comp_rfWrite <= Lsu2Plugin_logic_sq_mem_writeRd;
      end
      if(when_StateMachine_l253_1) begin
        Lsu2Plugin_logic_special_atomic_comp_wakeRf <= Lsu2Plugin_logic_sq_mem_writeRd;
        Lsu2Plugin_logic_special_atomic_comp_rfWrite <= (Lsu2Plugin_logic_special_storeSc && Lsu2Plugin_logic_sq_mem_writeRd);
      end
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_stateNext;
      if(DecoderPlugin_logic_exception_set) begin
        DecoderPlugin_logic_exception_trigged <= 1'b1;
      end
      if(DecoderPlugin_logic_exception_clear) begin
        DecoderPlugin_logic_exception_trigged <= 1'b0;
      end
      DecoderPlugin_logic_exception_doItAgain <= DecoderPlugin_logic_exception_doIt;
      FrontendPlugin_decoded_OP_ID <= (FrontendPlugin_decoded_OP_ID + _zz_FrontendPlugin_decoded_OP_ID);
      if(FrontendPlugin_serialized_valid) begin
        DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle <= 1'b0;
      end
      if(when_DecoderPredictionPlugin_l236) begin
        DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle <= 1'b1;
      end
      ALU0_ExecutionUnitBase_pipeline_fetch_1_valid <= ALU0_ExecutionUnitBase_pipeline_fetch_0_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        ALU0_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      end
      if(EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output) begin
        EU0_ExecutionUnitBase_pipeline_fetch_1_valid <= EU0_ExecutionUnitBase_pipeline_fetch_0_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        EU0_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      end
      if(EU0_ExecutionUnitBase_pipeline_execute_0_ready_output) begin
        EU0_ExecutionUnitBase_pipeline_execute_1_valid <= _zz_EU0_ExecutionUnitBase_pipeline_execute_1_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        EU0_ExecutionUnitBase_pipeline_execute_1_valid <= 1'b0;
      end
      if(EU0_ExecutionUnitBase_pipeline_execute_1_ready_output) begin
        EU0_ExecutionUnitBase_pipeline_execute_2_valid <= _zz_EU0_ExecutionUnitBase_pipeline_execute_2_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        EU0_ExecutionUnitBase_pipeline_execute_2_valid <= 1'b0;
      end
      if(BranchContextPlugin_free_learn_valid) begin
        BranchContextPlugin_logic_ptr_free <= (BranchContextPlugin_logic_ptr_free + 3'b001);
      end
      if(toplevel_DispatchPlugin_logic_queue_io_push_fire) begin
        DispatchPlugin_logic_ptr_next <= (DispatchPlugin_logic_ptr_next + 4'b0001);
        DispatchPlugin_logic_ptr_current <= (DispatchPlugin_logic_ptr_current + 4'b0001);
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        DispatchPlugin_logic_ptr_next <= (_zz_DispatchPlugin_logic_ptr_next + 4'b0001);
        DispatchPlugin_logic_ptr_current <= (CommitPlugin_logic_commit_reschedulePort_payload_robIdNext - 4'b1000);
      end
      if(when_DispatchPlugin_l192) begin
        DispatchPlugin_logic_push_fenceYoungerLast <= DispatchPlugin_logic_push_fenceYounger;
      end
      DispatchPlugin_logic_pop_0_stagesList_1_valid <= DispatchPlugin_logic_pop_0_stagesList_0_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        DispatchPlugin_logic_pop_0_stagesList_1_valid <= 1'b0;
      end
      if(DispatchPlugin_logic_pop_1_stagesList_0_ready_output) begin
        DispatchPlugin_logic_pop_1_stagesList_1_valid <= DispatchPlugin_logic_pop_1_stagesList_0_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        DispatchPlugin_logic_pop_1_stagesList_1_valid <= 1'b0;
      end
      if(RfDependencyPlugin_logic_forRf_integer_init_busy) begin
        RfDependencyPlugin_logic_forRf_integer_init_counter <= (RfDependencyPlugin_logic_forRf_integer_init_counter + 7'h01);
      end
      if(FrontendPlugin_allocated_ready_output) begin
        FrontendPlugin_dispatch_valid <= _zz_FrontendPlugin_dispatch_valid;
      end
      if(CommitPlugin_logic_reschedule_reschedulePort_valid) begin
        FrontendPlugin_dispatch_valid <= 1'b0;
      end
      if(FrontendPlugin_decoded_ready_output) begin
        FrontendPlugin_serialized_valid <= _zz_FrontendPlugin_serialized_valid;
      end
      if(when_Connection_l66) begin
        FrontendPlugin_serialized_valid <= 1'b0;
      end
      PcPlugin_logic_init_counter <= (PcPlugin_logic_init_counter + _zz_PcPlugin_logic_init_counter);
      if(PcPlugin_logic_fetchPc_correction) begin
        PcPlugin_logic_fetchPc_correctionReg <= 1'b1;
      end
      if(PcPlugin_logic_fetchPc_output_fire) begin
        PcPlugin_logic_fetchPc_correctionReg <= 1'b0;
      end
      if(when_PcPlugin_l84) begin
        PcPlugin_logic_fetchPc_inc <= 1'b0;
      end
      if(PcPlugin_logic_fetchPc_output_fire) begin
        PcPlugin_logic_fetchPc_inc <= 1'b1;
      end
      if(when_PcPlugin_l84_1) begin
        PcPlugin_logic_fetchPc_inc <= 1'b0;
      end
      if(when_PcPlugin_l100) begin
        PcPlugin_logic_fetchPc_pcReg <= PcPlugin_logic_fetchPc_pc;
      end
      if(when_Connection_l54) begin
        FetchPlugin_stages_1_valid <= 1'b0;
      end
      if(FetchPlugin_stages_0_ready_output) begin
        FetchPlugin_stages_1_valid <= _zz_FetchPlugin_stages_1_valid;
      end
      if(FetchPlugin_stages_1_ready_output) begin
        FetchPlugin_stages_2_valid <= _zz_FetchPlugin_stages_2_valid;
      end
      if(when_Connection_l66_1) begin
        FetchPlugin_stages_2_valid <= 1'b0;
      end
      if(_zz_AlignerPlugin_setup_s2m_valid) begin
        FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid <= 1'b1;
      end
      if(AlignerPlugin_setup_s2m_ready) begin
        FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid <= 1'b0;
      end
      if(FrontendPlugin_aligned_isFlushed) begin
        FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid <= 1'b0;
      end
      PrivilegedPlugin_logic_fsm_stateReg <= PrivilegedPlugin_logic_fsm_stateNext;
      case(PrivilegedPlugin_logic_fsm_stateReg)
        PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
          PrivilegedPlugin_setup_privilege <= PrivilegedPlugin_logic_fsm_xret_targetPrivilege;
          case(switch_PrivilegedPlugin_l960)
            2'b11 : begin
              PrivilegedPlugin_logic_machine_mstatus_mpp <= 2'b00;
              PrivilegedPlugin_logic_machine_mstatus_mie <= PrivilegedPlugin_logic_machine_mstatus_mpie;
              PrivilegedPlugin_logic_machine_mstatus_mpie <= 1'b1;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_supervisor_sstatus_spp <= 1'b0;
              PrivilegedPlugin_logic_supervisor_sstatus_sie <= PrivilegedPlugin_logic_supervisor_sstatus_spie;
              PrivilegedPlugin_logic_supervisor_sstatus_spie <= 1'b1;
            end
            default : begin
            end
          endcase
        end
        PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
          PrivilegedPlugin_setup_privilege <= PrivilegedPlugin_logic_fsm_trap_targetPrivilege;
          case(PrivilegedPlugin_logic_fsm_trap_targetPrivilege)
            2'b11 : begin
              PrivilegedPlugin_logic_machine_mstatus_mie <= 1'b0;
              PrivilegedPlugin_logic_machine_mstatus_mpie <= PrivilegedPlugin_logic_machine_mstatus_mie;
              PrivilegedPlugin_logic_machine_mstatus_mpp <= PrivilegedPlugin_setup_privilege;
              PrivilegedPlugin_logic_machine_cause_interrupt <= PrivilegedPlugin_logic_fsm_trap_interrupt;
              PrivilegedPlugin_logic_machine_cause_code <= PrivilegedPlugin_logic_fsm_trap_code;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_supervisor_sstatus_sie <= 1'b0;
              PrivilegedPlugin_logic_supervisor_sstatus_spie <= PrivilegedPlugin_logic_supervisor_sstatus_sie;
              PrivilegedPlugin_logic_supervisor_sstatus_spp <= PrivilegedPlugin_setup_privilege[0 : 0];
              PrivilegedPlugin_logic_supervisor_cause_interrupt <= PrivilegedPlugin_logic_fsm_trap_interrupt;
              PrivilegedPlugin_logic_supervisor_cause_code <= PrivilegedPlugin_logic_fsm_trap_code;
            end
            default : begin
            end
          endcase
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l253_2) begin
        PrivilegedPlugin_logic_decoderInterrupt_raised <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(when_FetchCachePlugin_l422) begin
      FetchCachePlugin_logic_refill_address <= FetchCachePlugin_logic_refill_start_address;
      FetchCachePlugin_logic_refill_isIo <= FetchCachePlugin_logic_refill_start_isIo;
    end
    if(AlignerPlugin_logic_fireInput) begin
      AlignerPlugin_logic_buffer_data <= AlignerPlugin_setup_s2m_Fetch_WORD;
      AlignerPlugin_logic_buffer_pc <= AlignerPlugin_setup_s2m_Fetch_FETCH_PC;
      AlignerPlugin_logic_buffer_fault <= AlignerPlugin_setup_s2m_Fetch_WORD_FAULT;
      AlignerPlugin_logic_buffer_fault_page <= AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE;
      AlignerPlugin_logic_buffer_branchValid <= (AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID && (! _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0));
      AlignerPlugin_logic_buffer_branchPcNext <= AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT;
      AlignerPlugin_logic_buffer_wordContexts_0 <= AlignerPlugin_setup_s2m_BRANCH_HISTORY;
      AlignerPlugin_logic_buffer_wordContexts_1 <= AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID;
      AlignerPlugin_logic_buffer_wordContexts_3 <= AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE;
      AlignerPlugin_logic_buffer_wordContexts_4_0 <= AlignerPlugin_setup_s2m_GSHARE_COUNTER_0;
      AlignerPlugin_logic_buffer_firstWordContexts_0 <= AlignerPlugin_setup_s2m_FETCH_ID;
    end
    CommitPlugin_logic_ptr_robLineMaskRsp <= CommitPlugin_setup_robLineMask_mask;
    if(when_CommitPlugin_l131) begin
      CommitPlugin_logic_reschedule_robId <= ((((_zz_CommitPlugin_logic_reschedule_trap ? Lsu2Plugin_setup_sharedTrap_payload_robId : 4'b0000) | (_zz_CommitPlugin_logic_reschedule_trap_1 ? Lsu2Plugin_setup_specialTrap_payload_robId : 4'b0000)) | ((_zz_CommitPlugin_logic_reschedule_trap_2 ? EU0_BranchPlugin_setup_reschedule_payload_robId : 4'b0000) | (_zz_CommitPlugin_logic_reschedule_trap_3 ? EnvCallPlugin_setup_reschedule_payload_robId : 4'b0000))) | (_zz_CommitPlugin_logic_reschedule_trap_4 ? EU0_CsrAccessPlugin_setup_trap_payload_robId : 4'b0000));
      CommitPlugin_logic_reschedule_trap <= _zz_CommitPlugin_logic_reschedule_trap_5[0];
      CommitPlugin_logic_reschedule_pcTarget <= ((CommitPlugin_logic_reschedule_portsLogic_hits[0] ? Lsu2Plugin_setup_sharedTrap_payload_pcTarget : 32'h00000000) | (CommitPlugin_logic_reschedule_portsLogic_hits[2] ? EU0_BranchPlugin_setup_reschedule_payload_pcTarget : 32'h00000000));
      CommitPlugin_logic_reschedule_cause <= ((((CommitPlugin_logic_reschedule_portsLogic_hits[0] ? Lsu2Plugin_setup_sharedTrap_payload_cause : 4'b0000) | (CommitPlugin_logic_reschedule_portsLogic_hits[1] ? Lsu2Plugin_setup_specialTrap_payload_cause : 4'b0000)) | ((CommitPlugin_logic_reschedule_portsLogic_hits[2] ? EU0_BranchPlugin_setup_reschedule_payload_cause : 4'b0000) | (CommitPlugin_logic_reschedule_portsLogic_hits[3] ? EnvCallPlugin_setup_reschedule_payload_cause : 4'b0000))) | (CommitPlugin_logic_reschedule_portsLogic_hits[4] ? EU0_CsrAccessPlugin_setup_trap_payload_cause : 4'b0000));
      CommitPlugin_logic_reschedule_reason <= ((((CommitPlugin_logic_reschedule_portsLogic_hits[0] ? Lsu2Plugin_setup_sharedTrap_payload_reason : 8'h00) | (CommitPlugin_logic_reschedule_portsLogic_hits[1] ? Lsu2Plugin_setup_specialTrap_payload_reason : 8'h00)) | ((CommitPlugin_logic_reschedule_portsLogic_hits[2] ? EU0_BranchPlugin_setup_reschedule_payload_reason : 8'h00) | (CommitPlugin_logic_reschedule_portsLogic_hits[3] ? EnvCallPlugin_setup_reschedule_payload_reason : 8'h00))) | (CommitPlugin_logic_reschedule_portsLogic_hits[4] ? EU0_CsrAccessPlugin_setup_trap_payload_reason : 8'h00));
      CommitPlugin_logic_reschedule_tval <= ((((CommitPlugin_logic_reschedule_portsLogic_hits[0] ? Lsu2Plugin_setup_sharedTrap_payload_tval : 32'h00000000) | (CommitPlugin_logic_reschedule_portsLogic_hits[1] ? Lsu2Plugin_setup_specialTrap_payload_tval : 32'h00000000)) | ((CommitPlugin_logic_reschedule_portsLogic_hits[2] ? EU0_BranchPlugin_setup_reschedule_payload_tval : 32'h00000000) | (CommitPlugin_logic_reschedule_portsLogic_hits[3] ? EnvCallPlugin_setup_reschedule_payload_tval : 32'h00000000))) | (CommitPlugin_logic_reschedule_portsLogic_hits[4] ? EU0_CsrAccessPlugin_setup_trap_payload_tval : 32'h00000000));
      CommitPlugin_logic_reschedule_skipCommit <= _zz_CommitPlugin_logic_reschedule_skipCommit[0];
    end
    PrivilegedPlugin_logic_supervisor_sip_seipInput <= PrivilegedPlugin_io_int_supervisor_external;
    if(PrivilegedPlugin_logic_rescheduleUnbuffered_ready) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_rData_cause <= PrivilegedPlugin_logic_rescheduleUnbuffered_payload_cause;
      PrivilegedPlugin_logic_rescheduleUnbuffered_rData_epc <= PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc;
      PrivilegedPlugin_logic_rescheduleUnbuffered_rData_tval <= PrivilegedPlugin_logic_rescheduleUnbuffered_payload_tval;
      PrivilegedPlugin_logic_rescheduleUnbuffered_rData_fromCommit <= PrivilegedPlugin_logic_rescheduleUnbuffered_payload_fromCommit;
    end
    if(LsuPlugin_peripheralBus_cmd_valid) begin
      LsuPlugin_peripheralBus_toAxiLite4_writeSel <= LsuPlugin_peripheralBus_cmd_payload_write;
    end
    if(DataCachePlugin_mem_toAxi4_awFiltred_ready) begin
      DataCachePlugin_mem_toAxi4_awFiltred_rData_last <= DataCachePlugin_mem_toAxi4_awFiltred_payload_last;
      DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_address <= DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_address;
      DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_data <= DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_data;
      DataCachePlugin_mem_toAxi4_awFiltred_rData_fragment_id <= DataCachePlugin_mem_toAxi4_awFiltred_payload_fragment_id;
    end
    if(Lsu2Plugin_logic_lq_regs_0_allocation) begin
      Lsu2Plugin_logic_lq_regs_0_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_1_allocation) begin
      Lsu2Plugin_logic_lq_regs_1_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_2_allocation) begin
      Lsu2Plugin_logic_lq_regs_2_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_3_allocation) begin
      Lsu2Plugin_logic_lq_regs_3_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_4_allocation) begin
      Lsu2Plugin_logic_lq_regs_4_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_5_allocation) begin
      Lsu2Plugin_logic_lq_regs_5_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_6_allocation) begin
      Lsu2Plugin_logic_lq_regs_6_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_7_allocation) begin
      Lsu2Plugin_logic_lq_regs_7_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_niceHazard <= 1'b0;
    end
    Lsu2Plugin_logic_lq_ptr_priorityLast <= Lsu2Plugin_logic_lq_ptr_priority;
    Lsu2Plugin_logic_lq_tracker_freeReduced <= _zz_Lsu2Plugin_logic_lq_tracker_freeReduced;
    if(Lsu2Plugin_logic_sq_regs_0_allocation) begin
      Lsu2Plugin_logic_sq_regs_0_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_1_allocation) begin
      Lsu2Plugin_logic_sq_regs_1_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_2_allocation) begin
      Lsu2Plugin_logic_sq_regs_2_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_3_allocation) begin
      Lsu2Plugin_logic_sq_regs_3_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_4_allocation) begin
      Lsu2Plugin_logic_sq_regs_4_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_5_allocation) begin
      Lsu2Plugin_logic_sq_regs_5_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_6_allocation) begin
      Lsu2Plugin_logic_sq_regs_6_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_7_allocation) begin
      Lsu2Plugin_logic_sq_regs_7_dataValid <= 1'b0;
    end
    Lsu2Plugin_logic_sq_ptr_priorityLast <= Lsu2Plugin_logic_sq_ptr_priority;
    Lsu2Plugin_logic_sq_ptr_onFreeLast_payload <= Lsu2Plugin_logic_sq_ptr_onFree_payload;
    Lsu2Plugin_logic_sq_tracker_freeReduced <= _zz_Lsu2Plugin_logic_sq_tracker_freeReduced;
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      case(switch_Utils_l1423)
        3'b000 : begin
          Lsu2Plugin_logic_lq_regs_0_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_0_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b001 : begin
          Lsu2Plugin_logic_lq_regs_1_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_1_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b010 : begin
          Lsu2Plugin_logic_lq_regs_2_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_2_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b011 : begin
          Lsu2Plugin_logic_lq_regs_3_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_3_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b100 : begin
          Lsu2Plugin_logic_lq_regs_4_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_4_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b101 : begin
          Lsu2Plugin_logic_lq_regs_5_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_5_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b110 : begin
          Lsu2Plugin_logic_lq_regs_6_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_6_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        default : begin
          Lsu2Plugin_logic_lq_regs_7_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_7_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
      endcase
    end
    if(when_Lsu2Plugin_l733) begin
      Lsu2Plugin_logic_sq_mem_swap <= AguPlugin_setup_port_payload_swap;
      Lsu2Plugin_logic_sq_mem_op <= AguPlugin_setup_port_payload_op;
      Lsu2Plugin_logic_sq_mem_physRd <= AguPlugin_setup_port_payload_physicalRd;
      Lsu2Plugin_logic_sq_mem_writeRd <= AguPlugin_setup_port_payload_writeRd;
    end
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      case(switch_Utils_l1423_1)
        3'b000 : begin
          Lsu2Plugin_logic_sq_regs_0_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_0_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_0_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b001 : begin
          Lsu2Plugin_logic_sq_regs_1_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_1_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_1_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b010 : begin
          Lsu2Plugin_logic_sq_regs_2_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_2_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_2_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b011 : begin
          Lsu2Plugin_logic_sq_regs_3_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_3_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_3_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b100 : begin
          Lsu2Plugin_logic_sq_regs_4_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_4_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_4_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b101 : begin
          Lsu2Plugin_logic_sq_regs_5_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_5_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_5_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        3'b110 : begin
          Lsu2Plugin_logic_sq_regs_6_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_6_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_6_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        default : begin
          Lsu2Plugin_logic_sq_regs_7_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_7_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_7_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
      endcase
    end
    if(when_Lsu2Plugin_l1046) begin
      case(Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID)
        3'b000 : begin
          Lsu2Plugin_logic_lq_regs_0_sqChecked <= 1'b1;
        end
        3'b001 : begin
          Lsu2Plugin_logic_lq_regs_1_sqChecked <= 1'b1;
        end
        3'b010 : begin
          Lsu2Plugin_logic_lq_regs_2_sqChecked <= 1'b1;
        end
        3'b011 : begin
          Lsu2Plugin_logic_lq_regs_3_sqChecked <= 1'b1;
        end
        3'b100 : begin
          Lsu2Plugin_logic_lq_regs_4_sqChecked <= 1'b1;
        end
        3'b101 : begin
          Lsu2Plugin_logic_lq_regs_5_sqChecked <= 1'b1;
        end
        3'b110 : begin
          Lsu2Plugin_logic_lq_regs_6_sqChecked <= 1'b1;
        end
        default : begin
          Lsu2Plugin_logic_lq_regs_7_sqChecked <= 1'b1;
        end
      endcase
    end
    if(when_Lsu2Plugin_l1104) begin
      Lsu2Plugin_logic_lq_regs_0_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_1) begin
      Lsu2Plugin_logic_lq_regs_1_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_2) begin
      Lsu2Plugin_logic_lq_regs_2_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_3) begin
      Lsu2Plugin_logic_lq_regs_3_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_4) begin
      Lsu2Plugin_logic_lq_regs_4_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_5) begin
      Lsu2Plugin_logic_lq_regs_5_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_6) begin
      Lsu2Plugin_logic_lq_regs_6_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_7) begin
      Lsu2Plugin_logic_lq_regs_7_niceHazard <= 1'b1;
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_118) begin
            Lsu2Plugin_logic_lq_regs_0_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_119) begin
            Lsu2Plugin_logic_lq_regs_1_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_120) begin
            Lsu2Plugin_logic_lq_regs_2_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_121) begin
            Lsu2Plugin_logic_lq_regs_3_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_122) begin
            Lsu2Plugin_logic_lq_regs_4_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_123) begin
            Lsu2Plugin_logic_lq_regs_5_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_124) begin
            Lsu2Plugin_logic_lq_regs_6_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_125) begin
            Lsu2Plugin_logic_lq_regs_7_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(when_Lsu2Plugin_l1333) begin
              if(Lsu2Plugin_logic_sharedPip_stages_3_LR) begin
                Lsu2Plugin_logic_lq_reservation_address <= Lsu2Plugin_logic_sharedPip_stages_3_MMU_TRANSLATED;
              end
            end
          end
        end
      endcase
    end
    if(Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready) begin
      toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rData <= Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_payload;
    end
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_fault <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_fault;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_redo <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_redo;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlot <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlot;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlotAny <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlotAny;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_generationKo <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_generationKo;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_flush <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_flush;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_prefetch <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_prefetch;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_address <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_address;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_io <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_io;
    if(Lsu2Plugin_setup_flushPort_cmd_valid) begin
      Lsu2Plugin_logic_flush_cmdPtr <= 3'b000;
      Lsu2Plugin_logic_flush_rspPtr <= 3'b000;
      Lsu2Plugin_logic_flush_withFree <= Lsu2Plugin_setup_flushPort_cmd_payload_withFree;
    end
    if(when_Lsu2Plugin_l1553) begin
      if(Lsu2Plugin_setup_cacheStore_cmd_fire) begin
        Lsu2Plugin_logic_flush_cmdPtr <= (Lsu2Plugin_logic_flush_cmdPtr + 3'b001);
      end
      if(when_Lsu2Plugin_l1561) begin
        if(Lsu2Plugin_setup_cacheStore_rsp_payload_redo) begin
          Lsu2Plugin_logic_flush_cmdPtr <= Lsu2Plugin_logic_flush_rspPtr;
        end else begin
          Lsu2Plugin_logic_flush_rspPtr <= (Lsu2Plugin_logic_flush_rspPtr + 3'b001);
        end
      end
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_isStore <= Lsu2Plugin_logic_special_storeHit;
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_isLoad <= (! Lsu2Plugin_logic_special_storeHit);
    end
    Lsu2Plugin_logic_special_robId <= CommitPlugin_logic_commit_head;
    Lsu2Plugin_logic_special_loadPhysRd <= Lsu2Plugin_logic_lq_mem_physRd_spinal_port2;
    Lsu2Plugin_logic_special_loadAddress <= Lsu2Plugin_logic_lq_mem_addressPost_spinal_port2;
    Lsu2Plugin_logic_special_loadAddressVirt <= Lsu2Plugin_logic_lq_mem_addressPre_spinal_port2;
    Lsu2Plugin_logic_special_loadSize <= Lsu2Plugin_logic_lq_mem_size_spinal_port2;
    Lsu2Plugin_logic_special_loadUnsigned <= Lsu2Plugin_logic_lq_mem_unsigned_spinal_port2[0];
    Lsu2Plugin_logic_special_loadWriteRd <= (Lsu2Plugin_logic_special_isLoad && Lsu2Plugin_logic_lq_mem_writeRd_spinal_port2[0]);
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeAddress <= Lsu2Plugin_setup_cacheStore_cmd_payload_address;
    end
    Lsu2Plugin_logic_special_storeAddressVirt <= Lsu2Plugin_logic_sq_mem_addressPre_spinal_port2;
    Lsu2Plugin_logic_special_storeSize <= Lsu2Plugin_logic_sq_mem_size_spinal_port4;
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeData <= Lsu2Plugin_setup_cacheStore_cmd_payload_data;
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeMask <= Lsu2Plugin_setup_cacheStore_cmd_payload_mask;
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeAmo <= Lsu2Plugin_logic_sq_mem_amo_spinal_port2[0];
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeSc <= Lsu2Plugin_logic_sq_mem_sc_spinal_port2[0];
    end
    if(PrivilegedPlugin_logic_decoderInterrupt_buffer_sample) begin
      PrivilegedPlugin_logic_decoderInterrupt_buffer_code <= PrivilegedPlugin_logic_interrupt_code;
    end
    if(PrivilegedPlugin_logic_decoderInterrupt_buffer_sample) begin
      PrivilegedPlugin_logic_decoderInterrupt_buffer_targetPrivilege <= PrivilegedPlugin_logic_interrupt_targetPrivilege;
    end
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
        EU0_CsrAccessPlugin_logic_fsm_regs_microOp <= EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
        EU0_CsrAccessPlugin_logic_fsm_regs_doImm <= EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_IMM;
        EU0_CsrAccessPlugin_logic_fsm_regs_doMask <= EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK;
        EU0_CsrAccessPlugin_logic_fsm_regs_doClear <= EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_CLEAR;
        EU0_CsrAccessPlugin_logic_fsm_regs_rs1 <= EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1;
        EU0_CsrAccessPlugin_logic_fsm_regs_implemented <= EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented;
        EU0_CsrAccessPlugin_logic_fsm_regs_trap <= EU0_CsrAccessPlugin_logic_fsm_startLogic_trap;
        EU0_CsrAccessPlugin_logic_fsm_regs_flushPipeline <= EU0_CsrAccessPlugin_setup_onDecodeFlushPipeline;
        EU0_CsrAccessPlugin_logic_fsm_regs_write <= EU0_CsrAccessPlugin_logic_fsm_startLogic_write;
        EU0_CsrAccessPlugin_logic_fsm_regs_read <= EU0_CsrAccessPlugin_logic_fsm_startLogic_read;
        REG_CSR_773 <= COMB_CSR_773;
        REG_CSR_835 <= COMB_CSR_835;
        REG_CSR_833 <= COMB_CSR_833;
        REG_CSR_832 <= COMB_CSR_832;
        REG_CSR_3857 <= COMB_CSR_3857;
        REG_CSR_3858 <= COMB_CSR_3858;
        REG_CSR_3859 <= COMB_CSR_3859;
        REG_CSR_3860 <= COMB_CSR_3860;
        REG_CSR_769 <= COMB_CSR_769;
        REG_CSR_834 <= COMB_CSR_834;
        REG_CSR_768 <= COMB_CSR_768;
        REG_CSR_836 <= COMB_CSR_836;
        REG_CSR_772 <= COMB_CSR_772;
        REG_CSR_770 <= COMB_CSR_770;
        REG_CSR_771 <= COMB_CSR_771;
        REG_CSR_261 <= COMB_CSR_261;
        REG_CSR_323 <= COMB_CSR_323;
        REG_CSR_321 <= COMB_CSR_321;
        REG_CSR_320 <= COMB_CSR_320;
        REG_CSR_322 <= COMB_CSR_322;
        REG_CSR_256 <= COMB_CSR_256;
        REG_CSR_260 <= COMB_CSR_260;
        REG_CSR_324 <= COMB_CSR_324;
        REG_CSR_384 <= COMB_CSR_384;
        EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b0;
        case(switch_CsrAccessPlugin_l206)
          12'h305 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 3'b111;
          end
          12'h343 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 3'b110;
          end
          12'h341 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 3'b101;
          end
          12'h340 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 3'b100;
          end
          12'h105 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 3'b011;
          end
          12'h143 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 3'b010;
          end
          12'h141 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 3'b001;
          end
          12'h140 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 3'b000;
          end
          default : begin
          end
        endcase
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        EU0_CsrAccessPlugin_logic_fsm_regs_aluInput <= EU0_CsrAccessPlugin_setup_onReadToWriteBits;
        EU0_CsrAccessPlugin_logic_fsm_regs_csrValue <= EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        if(EU0_CsrAccessPlugin_setup_onWriteFlushPipeline) begin
          EU0_CsrAccessPlugin_logic_fsm_regs_flushPipeline <= 1'b1;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
        if(EU0_ExecutionUnitBase_pipeline_execute_2_valid) begin
          EnvCallPlugin_logic_flushes_vmaInv <= EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA;
          EnvCallPlugin_logic_flushes_fetchInv <= EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I;
          EnvCallPlugin_logic_flushes_flushData <= EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
    MmuPlugin_logic_refill_portsOh_regNext <= MmuPlugin_logic_refill_portsOh;
    _zz_MmuPlugin_logic_refill_portsAddress <= Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION;
    _zz_MmuPlugin_logic_refill_portsAddress_1 <= FetchPlugin_stages_1_Fetch_FETCH_PC;
    MmuPlugin_logic_refill_load_rsp_payload_data <= MmuPlugin_setup_cacheLoad_rsp_payload_data;
    MmuPlugin_logic_refill_load_rsp_payload_fault <= MmuPlugin_setup_cacheLoad_rsp_payload_fault;
    MmuPlugin_logic_refill_load_rsp_payload_redo <= MmuPlugin_setup_cacheLoad_rsp_payload_redo;
    MmuPlugin_logic_refill_load_rsp_payload_refillSlot <= MmuPlugin_setup_cacheLoad_rsp_payload_refillSlot;
    MmuPlugin_logic_refill_load_rsp_payload_refillSlotAny <= MmuPlugin_setup_cacheLoad_rsp_payload_refillSlotAny;
    Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION <= Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION;
    Lsu2Plugin_logic_sharedPip_stages_1_ROB_ID <= Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_PHYS_RD <= Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD;
    Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_POST_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_1_SIZE <= Lsu2Plugin_logic_sharedPip_stages_0_SIZE;
    Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_1_TRANSLATED_AS_IO <= Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO;
    Lsu2Plugin_logic_sharedPip_stages_1_WRITE_RD <= Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD;
    Lsu2Plugin_logic_sharedPip_stages_1_UNSIGNED <= Lsu2Plugin_logic_sharedPip_stages_0_UNSIGNED;
    Lsu2Plugin_logic_sharedPip_stages_1_LR <= Lsu2Plugin_logic_sharedPip_stages_0_LR;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_VALID <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_DELTA <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SCORE <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SCORE;
    Lsu2Plugin_logic_sharedPip_stages_1_AMO <= Lsu2Plugin_logic_sharedPip_stages_0_AMO;
    Lsu2Plugin_logic_sharedPip_stages_1_SC <= Lsu2Plugin_logic_sharedPip_stages_0_SC;
    Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD <= Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD;
    Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID <= Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID <= Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH;
    Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION_COUNTER <= Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION_COUNTER;
    Lsu2Plugin_logic_sharedPip_stages_1_SP_FP_ADDRESS <= Lsu2Plugin_logic_sharedPip_stages_0_SP_FP_ADDRESS;
    Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK <= Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK;
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID <= Lsu2Plugin_logic_sharedPip_stages_0_LQCHECK_START_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID <= Lsu2Plugin_logic_sharedPip_stages_0_SQCHECK_END_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE <= Lsu2Plugin_logic_sharedPip_stages_0_feed_SQ_PTR_FREE;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SQID <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SQID;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_FEEDED;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH_PC <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH_PC;
    Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL <= Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL_overloaded;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS_PRE_VALID <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_HITS_PRE_VALID;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SQID <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SQID;
    Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_TRANSLATED <= Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED;
    Lsu2Plugin_logic_sharedPip_stages_2_IS_IO <= Lsu2Plugin_logic_sharedPip_stages_1_IS_IO;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_TRANSLATED <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_ACCESS_FAULT <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_READ <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_REDO <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO;
    Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_HIT <= Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_HIT;
    Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID <= Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_ID;
    Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD <= Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT;
    Lsu2Plugin_logic_sharedPip_stages_2_LQ_ID <= Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_2_SQ_ID <= Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS <= Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS;
    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_NO_YOUNGER <= Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_WRITE <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_WRITE;
    Lsu2Plugin_logic_sharedPip_stages_2_SIZE <= Lsu2Plugin_logic_sharedPip_stages_1_SIZE;
    Lsu2Plugin_logic_sharedPip_stages_2_UNSIGNED <= Lsu2Plugin_logic_sharedPip_stages_1_UNSIGNED;
    Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID <= Lsu2Plugin_logic_sharedPip_stages_1_ROB_ID;
    Lsu2Plugin_logic_sharedPip_stages_2_WRITE_RD <= Lsu2Plugin_logic_sharedPip_stages_1_WRITE_RD;
    Lsu2Plugin_logic_sharedPip_stages_2_PHYS_RD <= Lsu2Plugin_logic_sharedPip_stages_1_PHYS_RD;
    Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION <= Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION;
    Lsu2Plugin_logic_sharedPip_stages_2_LR <= Lsu2Plugin_logic_sharedPip_stages_1_LR;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SCORE <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SCORE;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_VALID <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_VALID;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_DELTA <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_DELTA;
    Lsu2Plugin_logic_sharedPip_stages_2_SC <= Lsu2Plugin_logic_sharedPip_stages_1_SC;
    Lsu2Plugin_logic_sharedPip_stages_2_AMO <= Lsu2Plugin_logic_sharedPip_stages_1_AMO;
    Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION_COUNTER <= Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION_COUNTER;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH;
    Lsu2Plugin_logic_sharedPip_stages_2_SP_FP_ADDRESS <= Lsu2Plugin_logic_sharedPip_stages_1_SP_FP_ADDRESS;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH_PC <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH_PC;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SQID <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SQID;
    Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED <= Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED_overloaded;
    Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID <= Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_WAIT_FEED <= Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED;
    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ROB <= Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ROB;
    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE <= Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_RESCHEDULE;
    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ID <= Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_valid <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_valid;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_data <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_data;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_fault <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_fault;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_redo <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_redo;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlot <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlot;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlotAny <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny;
    Lsu2Plugin_logic_sharedPip_stages_3_ADDRESS_PRE_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_3_IS_IO <= Lsu2Plugin_logic_sharedPip_stages_2_IS_IO;
    Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD <= Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD;
    Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID <= Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID <= Lsu2Plugin_logic_sharedPip_stages_2_LQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_WRITE_RD <= Lsu2Plugin_logic_sharedPip_stages_2_WRITE_RD;
    Lsu2Plugin_logic_sharedPip_stages_3_PHYS_RD <= Lsu2Plugin_logic_sharedPip_stages_2_PHYS_RD;
    Lsu2Plugin_logic_sharedPip_stages_3_CTRL <= Lsu2Plugin_logic_sharedPip_stages_2_CTRL;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT;
    Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION <= Lsu2Plugin_logic_sharedPip_stages_2_TRAP_SPECULATION;
    Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION <= Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION;
    Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID <= Lsu2Plugin_logic_sharedPip_stages_2_SQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_LR <= Lsu2Plugin_logic_sharedPip_stages_2_LR;
    Lsu2Plugin_logic_sharedPip_stages_3_MMU_TRANSLATED <= Lsu2Plugin_logic_sharedPip_stages_2_MMU_TRANSLATED;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SCORE;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_VALID <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_VALID;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_DELTA <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_DELTA;
    Lsu2Plugin_logic_sharedPip_stages_3_SC <= Lsu2Plugin_logic_sharedPip_stages_2_SC;
    Lsu2Plugin_logic_sharedPip_stages_3_AMO <= Lsu2Plugin_logic_sharedPip_stages_2_AMO;
    Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION_COUNTER <= Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION_COUNTER;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH;
    Lsu2Plugin_logic_sharedPip_stages_3_SP_FP_ADDRESS <= Lsu2Plugin_logic_sharedPip_stages_2_SP_FP_ADDRESS;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH_PC <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH_PC;
    if(Lsu2Plugin_logic_lqSqArbitration_s0_ready_output) begin
      Lsu2Plugin_logic_lqSqArbitration_s1_LQ_HIT <= Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT;
      Lsu2Plugin_logic_lqSqArbitration_s1_SQ_HIT <= Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT;
      Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID <= Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID;
      Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID <= Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID;
      Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ROB_FULL <= Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ROB_FULL;
      Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ROB_FULL <= Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ROB_FULL;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_IDLE_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP_OH_ID]) : begin
        Lsu2Plugin_logic_special_atomic_readed <= Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated[31 : 0];
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY_OH_ID]) : begin
        if(when_Lsu2Plugin_l1715) begin
          Lsu2Plugin_logic_special_atomic_gotReservation <= (Lsu2Plugin_logic_lq_reservation_valid && (Lsu2Plugin_logic_lq_reservation_address == Lsu2Plugin_logic_special_storeAddress));
        end
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_ALU_OH_ID]) : begin
        Lsu2Plugin_logic_special_atomic_result <= Lsu2Plugin_logic_special_atomic_alu_result;
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_SYNC_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_OH_ID]) : begin
      end
      (Lsu2Plugin_logic_special_atomic_stateReg[Lsu2Plugin_logic_special_atomic_enumDef_TRAP_WAIT_OH_ID]) : begin
      end
      default : begin
      end
    endcase
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
        MmuPlugin_logic_refill_portOhReg <= MmuPlugin_logic_refill_portsOh;
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
        MmuPlugin_logic_refill_virtual <= MmuPlugin_logic_refill_portsAddress;
        MmuPlugin_logic_refill_load_address <= {{MmuPlugin_logic_satp_ppn,MmuPlugin_logic_refill_portsAddress[31 : 22]},2'b00};
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(!when_MmuPlugin_l499) begin
              MmuPlugin_logic_refill_load_address <= MmuPlugin_logic_refill_load_nextLevelBase;
              MmuPlugin_logic_refill_load_address[11 : 2] <= MmuPlugin_logic_refill_virtual[21 : 12];
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(when_DecoderPlugin_l302) begin
      DecoderPlugin_logic_exception_exceptionReg_0 <= FrontendPlugin_decoded_TRAP_0;
    end
    if(when_DecoderPlugin_l303) begin
      DecoderPlugin_logic_exception_fetchFaultReg_0 <= FrontendPlugin_decoded_Frontend_FETCH_FAULT_0;
    end
    if(when_DecoderPlugin_l304) begin
      DecoderPlugin_logic_exception_fetchFaultPageReg_0 <= FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_0;
    end
    if(when_DecoderPlugin_l306) begin
      DecoderPlugin_logic_exception_debugEnterReg_0 <= DecoderPlugin_setup_debugEnter_0;
    end
    if(when_DecoderPlugin_l307) begin
      DecoderPlugin_logic_exception_epcReg_0 <= FrontendPlugin_decoded_PC_0;
    end
    if(when_DecoderPlugin_l308) begin
      DecoderPlugin_logic_exception_instReg_0 <= FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_0;
    end
    if(when_DecoderPlugin_l309) begin
      DecoderPlugin_logic_exception_compressedFaultReg_0 <= FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_0;
    end
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1 <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2 <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID <= ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD <= ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD <= ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0 <= ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT <= ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED <= ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
    if(EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output) begin
      EU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP <= EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1 <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
      EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS1 <= EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2 <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
      EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS2 <= EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
      EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID <= EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
      EU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD <= EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
      EU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD <= EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
      EU0_ExecutionUnitBase_pipeline_fetch_1_PC <= EU0_ExecutionUnitBase_pipeline_fetch_0_PC;
      EU0_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID <= EU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
      EU0_ExecutionUnitBase_pipeline_fetch_1_LSU_ID <= EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID;
      EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_MSB <= EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB;
      EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E2 <= EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2;
      EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_HIGH <= EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH;
      EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS1_SIGNED <= EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED;
      EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS2_SIGNED <= EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED;
      EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_REM <= EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM;
      EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL <= EU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_AMO <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SC <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LOAD <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LR <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_ECALL <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_EBREAK <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_XRET <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_WFI <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_I <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_VMA <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FLUSH_DATA <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA;
      EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_IMM <= EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM;
      EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_MASK <= EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK;
      EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_CLEAR <= EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_0_ready_output) begin
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_0;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_1;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_2 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_2;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_3 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_3;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_4 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_4;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_5 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_5;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_6 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_6;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_7 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_7;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_8 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_8;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_9 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_9;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_10 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_10;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_11 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_11;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_12 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_12;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_13 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_13;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_14 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_14;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_15 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_15;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_16 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_16;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_17 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_17;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_18 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_18;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_19 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_19;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_20 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_20;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_21 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_21;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_22 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_22;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_23 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_23;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_24 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_24;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_25 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_25;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_26 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_26;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_27 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_27;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_28 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_28;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_29 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_29;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_30 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_30;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_31 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_31;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_32 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_32;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_33 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_33;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_34 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_34;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_35 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_35;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_36 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_36;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_37 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_37;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_38 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_38;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_39 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_39;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_40 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_40;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_41 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_41;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_42 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_42;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_43 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_43;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_44 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_44;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_45 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_45;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_46 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_46;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_47 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_47;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_48 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_48;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_49 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_49;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_50 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_50;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_51 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_51;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_52 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_52;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_53 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_53;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_54 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_54;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_55 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_55;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_56 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_56;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_57 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_57;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_58 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_58;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_59 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_59;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_60 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_60;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_61 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_61;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_62 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_62;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_63 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_63;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_64 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_64;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_65 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_steps_0_adders_65;
      EU0_ExecutionUnitBase_pipeline_execute_1_DIV_REVERT_RESULT <= EU0_ExecutionUnitBase_pipeline_execute_0_DIV_REVERT_RESULT;
      EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_REM <= EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM;
      EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND <= EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
      EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL <= EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL;
      EU0_ExecutionUnitBase_pipeline_execute_1_Frontend_MICRO_OP <= EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
      EU0_ExecutionUnitBase_pipeline_execute_1_PC <= EU0_ExecutionUnitBase_pipeline_execute_0_PC;
      EU0_ExecutionUnitBase_pipeline_execute_1_PC_TRUE <= EU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
      EU0_ExecutionUnitBase_pipeline_execute_1_PC_FALSE <= EU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE;
      EU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET <= EU0_ExecutionUnitBase_pipeline_execute_0_PC_TARGET;
      EU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken <= EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
      EU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_pc <= EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc;
      EU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID <= EU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID;
      EU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID <= EU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
      EU0_ExecutionUnitBase_pipeline_execute_1_PHYS_RD <= EU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
      EU0_ExecutionUnitBase_pipeline_execute_1_WRITE_RD <= EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
      EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET <= EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET;
      EU0_ExecutionUnitBase_pipeline_execute_1_CsrAccessPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_HIGH <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_HIGH;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_EBREAK <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_EBREAK;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_ECALL <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_ECALL;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_XRET <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_XRET;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_I <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_I;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FLUSH_DATA <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FLUSH_DATA;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_VMA <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_VMA;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_WFI <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_WFI;
      EU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E2 <= EU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E2;
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_1_ready_output) begin
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_0;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_1 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_1;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_2 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_2;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_3 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_3;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_4 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_4;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_5 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_5;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_6 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_6;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_7 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_7;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_8 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_8;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_9 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_1_adders_9;
      EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_DIV_RESULT <= EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT;
      EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID <= EU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
      EU0_ExecutionUnitBase_pipeline_execute_2_BranchPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_2_PC <= EU0_ExecutionUnitBase_pipeline_execute_1_PC;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_HIGH <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_HIGH;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_EBREAK;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_ECALL;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_XRET;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_I;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FLUSH_DATA;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_VMA;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_WFI <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_WFI;
      EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_1_CsrAccessPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_2_PC_FALSE <= EU0_ExecutionUnitBase_pipeline_execute_1_PC_FALSE;
      EU0_ExecutionUnitBase_pipeline_execute_2_Frontend_MICRO_OP <= EU0_ExecutionUnitBase_pipeline_execute_1_Frontend_MICRO_OP;
      EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD <= EU0_ExecutionUnitBase_pipeline_execute_1_WRITE_RD;
      EU0_ExecutionUnitBase_pipeline_execute_2_PHYS_RD <= EU0_ExecutionUnitBase_pipeline_execute_1_PHYS_RD;
      EU0_ExecutionUnitBase_pipeline_execute_2_completion_SEL_E2 <= EU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E2;
    end
    DispatchPlugin_logic_pop_0_stagesList_1_OFFSET <= DispatchPlugin_logic_pop_0_stagesList_0_OFFSET;
    DispatchPlugin_logic_pop_0_stagesList_1_UINT <= DispatchPlugin_logic_pop_0_stagesList_0_UINT;
    DispatchPlugin_logic_pop_0_stagesList_1_LATENCY_0 <= DispatchPlugin_logic_pop_0_stagesList_0_LATENCY_0;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_0 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_1 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_2 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_3 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3;
    if(DispatchPlugin_logic_pop_1_stagesList_0_ready_output) begin
      DispatchPlugin_logic_pop_1_stagesList_1_OFFSET <= DispatchPlugin_logic_pop_1_stagesList_0_OFFSET;
      DispatchPlugin_logic_pop_1_stagesList_1_UINT <= DispatchPlugin_logic_pop_1_stagesList_0_UINT;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_0 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_0;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_1 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_1;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_2 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_2;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RD_3 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RD_3;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_0 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_0;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_1 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_1;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_2 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_2;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_0_3 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_0_3;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_0 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_0;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_1 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_1;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_2 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_2;
      DispatchPlugin_logic_pop_1_stagesList_1_EU0_readContext_PHYS_RS_1_3 <= DispatchPlugin_logic_pop_1_stagesList_0_EU0_readContext_PHYS_RS_1_3;
    end
    if(FrontendPlugin_allocated_ready_output) begin
      FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 <= FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0;
      FrontendPlugin_dispatch_WRITE_RD_0 <= FrontendPlugin_allocated_WRITE_RD_0;
      FrontendPlugin_dispatch_PHYS_RD_0 <= FrontendPlugin_allocated_PHYS_RD_0;
      FrontendPlugin_dispatch_BRANCH_ID_0 <= FrontendPlugin_allocated_BRANCH_ID_0;
      FrontendPlugin_dispatch_BRANCH_SEL_0 <= FrontendPlugin_allocated_BRANCH_SEL_0;
      FrontendPlugin_dispatch_ROB_ID <= FrontendPlugin_allocated_ROB_ID;
      FrontendPlugin_dispatch_ARCH_RS_0_0 <= FrontendPlugin_allocated_ARCH_RS_0_0;
      FrontendPlugin_dispatch_READ_RS_0_0 <= FrontendPlugin_allocated_READ_RS_0_0;
      FrontendPlugin_dispatch_PHYS_RS_0_0 <= FrontendPlugin_allocated_PHYS_RS_0_0;
      FrontendPlugin_dispatch_READ_RS_1_0 <= FrontendPlugin_allocated_READ_RS_1_0;
      FrontendPlugin_dispatch_PHYS_RS_1_0 <= FrontendPlugin_allocated_PHYS_RS_1_0;
      FrontendPlugin_dispatch_BRANCH_HISTORY_0 <= FrontendPlugin_allocated_BRANCH_HISTORY_0;
      FrontendPlugin_dispatch_Frontend_MICRO_OP_0 <= FrontendPlugin_allocated_Frontend_MICRO_OP_0;
      FrontendPlugin_dispatch_LQ_ALLOC_0 <= FrontendPlugin_allocated_LQ_ALLOC_0;
      FrontendPlugin_dispatch_SQ_ALLOC_0 <= FrontendPlugin_allocated_SQ_ALLOC_0;
      FrontendPlugin_dispatch_Prediction_IS_BRANCH_0 <= FrontendPlugin_allocated_Prediction_IS_BRANCH_0;
      FrontendPlugin_dispatch_GSHARE_COUNTER_0_0 <= FrontendPlugin_allocated_GSHARE_COUNTER_0_0;
      FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_0 <= FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_0;
      FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_0 <= FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_0;
      FrontendPlugin_dispatch_ALU0_SEL_0 <= FrontendPlugin_allocated_ALU0_SEL_0;
      FrontendPlugin_dispatch_EU0_SEL_0 <= FrontendPlugin_allocated_EU0_SEL_0;
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_0 <= FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_0;
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_0 <= FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_0;
    end
    if(FrontendPlugin_decoded_ready_output) begin
      FrontendPlugin_serialized_FETCH_ID_0 <= FrontendPlugin_decoded_FETCH_ID_0;
      FrontendPlugin_serialized_READ_RS_0_0 <= FrontendPlugin_decoded_READ_RS_0_0;
      FrontendPlugin_serialized_READ_RS_1_0 <= FrontendPlugin_decoded_READ_RS_1_0;
      FrontendPlugin_serialized_WRITE_RD_0 <= FrontendPlugin_decoded_WRITE_RD_0;
      FrontendPlugin_serialized_ALU0_SEL_0 <= FrontendPlugin_decoded_ALU0_SEL_0;
      FrontendPlugin_serialized_EU0_SEL_0 <= FrontendPlugin_decoded_EU0_SEL_0;
      FrontendPlugin_serialized_LQ_ALLOC_0 <= FrontendPlugin_decoded_LQ_ALLOC_0;
      FrontendPlugin_serialized_SQ_ALLOC_0 <= FrontendPlugin_decoded_SQ_ALLOC_0;
      FrontendPlugin_serialized_Frontend_DECODED_MASK_0 <= FrontendPlugin_decoded_Frontend_DECODED_MASK_0;
      FrontendPlugin_serialized_Frontend_MICRO_OP_0 <= FrontendPlugin_decoded_Frontend_MICRO_OP_0;
      FrontendPlugin_serialized_ARCH_RD_0 <= FrontendPlugin_decoded_ARCH_RD_0;
      FrontendPlugin_serialized_ARCH_RS_0_0 <= FrontendPlugin_decoded_ARCH_RS_0_0;
      FrontendPlugin_serialized_ARCH_RS_1_0 <= FrontendPlugin_decoded_ARCH_RS_1_0;
      FrontendPlugin_serialized_PC_0 <= FrontendPlugin_decoded_PC_0;
      FrontendPlugin_serialized_OP_ID <= FrontendPlugin_decoded_OP_ID;
      FrontendPlugin_serialized_IS_JALR_0 <= FrontendPlugin_decoded_IS_JALR_0;
      FrontendPlugin_serialized_Prediction_IS_BRANCH_0 <= FrontendPlugin_decoded_Prediction_IS_BRANCH_0;
      FrontendPlugin_serialized_IS_ANY_0 <= FrontendPlugin_decoded_IS_ANY_0;
      FrontendPlugin_serialized_RAS_PUSH_0 <= FrontendPlugin_decoded_RAS_PUSH_0;
      FrontendPlugin_serialized_RAS_POP_0 <= FrontendPlugin_decoded_RAS_POP_0;
      FrontendPlugin_serialized_PC_INC_0 <= FrontendPlugin_decoded_PC_INC_0;
      FrontendPlugin_serialized_PC_TARGET_PRE_RAS_0 <= FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0;
      FrontendPlugin_serialized_BAD_RET_PC_0 <= FrontendPlugin_decoded_BAD_RET_PC_0;
      FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_0 <= FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
      FrontendPlugin_serialized_CAN_IMPROVE_0 <= FrontendPlugin_decoded_CAN_IMPROVE_0;
      FrontendPlugin_serialized_BRANCHED_PREDICTION_0 <= FrontendPlugin_decoded_BRANCHED_PREDICTION_0;
      FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0 <= FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_0;
      FrontendPlugin_serialized_BRANCH_HISTORY_0 <= FrontendPlugin_decoded_BRANCH_HISTORY_0;
      FrontendPlugin_serialized_GSHARE_COUNTER_0_0 <= FrontendPlugin_decoded_GSHARE_COUNTER_0_0;
    end
    if(FetchPlugin_stages_0_ready_output) begin
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_loaded <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_error <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_error;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_address;
      FetchPlugin_stages_1_Fetch_FETCH_PC <= FetchPlugin_stages_0_Fetch_FETCH_PC;
      FetchPlugin_stages_1_GSharePlugin_logic_HASH <= FetchPlugin_stages_0_GSharePlugin_logic_HASH;
      FetchPlugin_stages_1_BRANCH_HISTORY <= FetchPlugin_stages_0_BRANCH_HISTORY;
      FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_valid <= FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_valid;
      FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_address <= FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_address;
      FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_0 <= FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_0;
    end
    if(FetchPlugin_stages_1_ready_output) begin
      FetchPlugin_stages_2_FETCH_ID <= FetchPlugin_stages_1_FETCH_ID;
      FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_0 <= FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_0;
      FetchPlugin_stages_2_Fetch_FETCH_PC <= FetchPlugin_stages_1_Fetch_FETCH_PC;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_loaded <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_error <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_error;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_address <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_0 <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_0;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HIT <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HIT;
      FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT <= FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT;
      FetchPlugin_stages_2_GSHARE_COUNTER_0 <= FetchPlugin_stages_1_GSHARE_COUNTER_0;
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID <= FetchPlugin_stages_1_Prediction_WORD_BRANCH_VALID;
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT <= FetchPlugin_stages_1_Prediction_WORD_BRANCH_PC_NEXT;
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID <= FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALID;
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE <= FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALUE;
      FetchPlugin_stages_2_MMU_IO <= FetchPlugin_stages_1_MMU_IO;
      FetchPlugin_stages_2_MMU_TRANSLATED <= FetchPlugin_stages_1_MMU_TRANSLATED;
      FetchPlugin_stages_2_MMU_REDO <= FetchPlugin_stages_1_MMU_REDO;
      FetchPlugin_stages_2_MMU_ALLOW_EXECUTE <= FetchPlugin_stages_1_MMU_ALLOW_EXECUTE;
      FetchPlugin_stages_2_MMU_PAGE_FAULT <= FetchPlugin_stages_1_MMU_PAGE_FAULT;
      FetchPlugin_stages_2_MMU_ACCESS_FAULT <= FetchPlugin_stages_1_MMU_ACCESS_FAULT;
      FetchPlugin_stages_2_Fetch_FETCH_PC_INC <= FetchPlugin_stages_1_Fetch_FETCH_PC_INC;
      FetchPlugin_stages_2_BRANCH_HISTORY <= FetchPlugin_stages_1_BRANCH_HISTORY;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_WORD_s2mBuffer <= FetchPlugin_stages_2_Fetch_WORD;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_FETCH_PC_s2mBuffer <= FetchPlugin_stages_2_Fetch_FETCH_PC;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_WORD_FAULT_s2mBuffer <= FetchPlugin_stages_2_Fetch_WORD_FAULT;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE_s2mBuffer <= FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_BRANCH_HISTORY_s2mBuffer <= FetchPlugin_stages_2_BRANCH_HISTORY;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_FETCH_ID_s2mBuffer <= FetchPlugin_stages_2_FETCH_ID;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID_s2mBuffer <= FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT_s2mBuffer <= FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT_s2mBuffer <= FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID_s2mBuffer <= FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE_s2mBuffer <= FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_0 <= FetchPlugin_stages_2_GSHARE_COUNTER_0;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_FETCH_PC_INC_s2mBuffer <= FetchPlugin_stages_2_Fetch_FETCH_PC_INC;
    end
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
        if(when_PrivilegedPlugin_l773) begin
          PrivilegedPlugin_logic_fsm_trap_interrupt <= 1'b1;
          PrivilegedPlugin_logic_fsm_trap_code <= PrivilegedPlugin_logic_decoderInterrupt_buffer_code;
          PrivilegedPlugin_logic_fsm_trap_targetPrivilege <= PrivilegedPlugin_logic_decoderInterrupt_buffer_targetPrivilege;
        end else begin
          case(PrivilegedPlugin_logic_reschedule_payload_cause)
            4'b1001 : begin
            end
            4'b1010 : begin
            end
            4'b1000 : begin
            end
            default : begin
              PrivilegedPlugin_logic_fsm_trap_interrupt <= 1'b0;
              PrivilegedPlugin_logic_fsm_trap_code <= PrivilegedPlugin_logic_exception_code;
              PrivilegedPlugin_logic_fsm_trap_targetPrivilege <= PrivilegedPlugin_logic_exception_targetPrivilege;
            end
          endcase
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        PrivilegedPlugin_logic_readed <= PrivilegedPlugin_setup_ramRead_data;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        PrivilegedPlugin_logic_readed <= PrivilegedPlugin_setup_ramRead_data;
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
        PrivilegedPlugin_logic_readed[31 : 0] <= _zz_PrivilegedPlugin_logic_readed;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end


endmodule

module DependencyStorage (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_payload_physical,
  input  wire [3:0]    io_writes_0_payload_robId,
  input  wire          io_commits_0_valid,
  input  wire [5:0]    io_commits_0_payload_physical,
  input  wire          io_commits_1_valid,
  input  wire [5:0]    io_commits_1_payload_physical,
  input  wire          io_commits_2_valid,
  input  wire [5:0]    io_commits_2_payload_physical,
  input  wire          io_commits_3_valid,
  input  wire [5:0]    io_commits_3_payload_physical,
  input  wire          io_commits_4_valid,
  input  wire [5:0]    io_commits_4_payload_physical,
  input  wire          io_reads_0_cmd_valid,
  input  wire [5:0]    io_reads_0_cmd_payload,
  output wire          io_reads_0_rsp_valid,
  output wire          io_reads_0_rsp_payload_enable,
  output wire [3:0]    io_reads_0_rsp_payload_rob,
  input  wire          io_reads_1_cmd_valid,
  input  wire [5:0]    io_reads_1_cmd_payload,
  output wire          io_reads_1_rsp_valid,
  output wire          io_reads_1_rsp_payload_enable,
  output wire [3:0]    io_reads_1_rsp_payload_rob,
  input  wire          clk,
  input  wire          reset
);

  wire       [3:0]    translation_physToRob_spinal_port1;
  wire       [3:0]    translation_physToRob_spinal_port2;
  wire       [3:0]    _zz_translation_physToRob_port;
  wire       [63:0]   _zz_status_sets;
  wire       [63:0]   _zz_status_clears;
  wire       [63:0]   _zz_status_clears_1;
  wire       [63:0]   _zz_status_clears_2;
  wire       [63:0]   _zz_status_clears_3;
  wire       [63:0]   _zz_status_clears_4;
  reg        [63:0]   status_busy;
  wire       [63:0]   status_sets;
  wire       [63:0]   status_clears;
  wire       [3:0]    read_0_robId;
  wire                read_0_enabled;
  wire       [3:0]    read_1_robId;
  wire                read_1_enabled;
  (* ram_style = "distributed" *) reg [3:0] translation_physToRob [0:63];

  assign _zz_status_sets = (64'h0000000000000001 <<< io_writes_0_payload_physical);
  assign _zz_status_clears = (64'h0000000000000001 <<< io_commits_0_payload_physical);
  assign _zz_status_clears_1 = (64'h0000000000000001 <<< io_commits_1_payload_physical);
  assign _zz_status_clears_2 = (64'h0000000000000001 <<< io_commits_2_payload_physical);
  assign _zz_status_clears_3 = (64'h0000000000000001 <<< io_commits_3_payload_physical);
  assign _zz_status_clears_4 = (64'h0000000000000001 <<< io_commits_4_payload_physical);
  assign _zz_translation_physToRob_port = io_writes_0_payload_robId;
  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      translation_physToRob[io_writes_0_payload_physical] <= _zz_translation_physToRob_port;
    end
  end

  assign translation_physToRob_spinal_port1 = translation_physToRob[io_reads_0_cmd_payload];
  assign translation_physToRob_spinal_port2 = translation_physToRob[io_reads_1_cmd_payload];
  assign status_sets = (io_writes_0_valid ? _zz_status_sets : 64'h0000000000000000);
  assign status_clears = ((((io_commits_0_valid ? _zz_status_clears : 64'h0000000000000000) | (io_commits_1_valid ? _zz_status_clears_1 : 64'h0000000000000000)) | ((io_commits_2_valid ? _zz_status_clears_2 : 64'h0000000000000000) | (io_commits_3_valid ? _zz_status_clears_3 : 64'h0000000000000000))) | (io_commits_4_valid ? _zz_status_clears_4 : 64'h0000000000000000));
  assign read_0_robId = translation_physToRob_spinal_port1;
  assign read_0_enabled = status_busy[io_reads_0_cmd_payload];
  assign io_reads_0_rsp_valid = io_reads_0_cmd_valid;
  assign io_reads_0_rsp_payload_enable = read_0_enabled;
  assign io_reads_0_rsp_payload_rob = read_0_robId;
  assign read_1_robId = translation_physToRob_spinal_port2;
  assign read_1_enabled = status_busy[io_reads_1_cmd_payload];
  assign io_reads_1_rsp_valid = io_reads_1_cmd_valid;
  assign io_reads_1_rsp_payload_enable = read_1_enabled;
  assign io_reads_1_rsp_payload_rob = read_1_robId;
  always @(posedge clk) begin
    status_busy <= ((status_busy & (~ status_clears)) | status_sets);
  end


endmodule

module RegFileLatch (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_address,
  input  wire [31:0]   io_writes_0_data,
  input  wire [3:0]    io_writes_0_robId,
  input  wire          io_writes_1_valid,
  input  wire [5:0]    io_writes_1_address,
  input  wire [31:0]   io_writes_1_data,
  input  wire [3:0]    io_writes_1_robId,
  input  wire          io_reads_0_valid,
  input  wire [5:0]    io_reads_0_address,
  output wire [31:0]   io_reads_0_data,
  input  wire          io_reads_1_valid,
  input  wire [5:0]    io_reads_1_address,
  output wire [31:0]   io_reads_1_data,
  input  wire          io_reads_2_valid,
  input  wire [5:0]    io_reads_2_address,
  output wire [31:0]   io_reads_2_data,
  input  wire          io_reads_3_valid,
  input  wire [5:0]    io_reads_3_address,
  output wire [31:0]   io_reads_3_data,
  input  wire          clk,
  input  wire          reset
);

  wire       [31:0]   _zz_readLogic_0_tri_64;
  wire       [31:0]   _zz_readLogic_1_tri_64;
  wire       [31:0]   _zz_readLogic_2_tri_64;
  wire       [31:0]   _zz_readLogic_3_tri_64;
  reg                 _zz_readLogic_3_tri;
  reg                 _zz_readLogic_3_tri_1;
  reg                 _zz_readLogic_3_tri_2;
  reg                 _zz_readLogic_3_tri_3;
  reg                 _zz_readLogic_3_tri_4;
  reg                 _zz_readLogic_3_tri_5;
  reg                 _zz_readLogic_3_tri_6;
  reg                 _zz_readLogic_3_tri_7;
  reg                 _zz_readLogic_3_tri_8;
  reg                 _zz_readLogic_3_tri_9;
  reg                 _zz_readLogic_3_tri_10;
  reg                 _zz_readLogic_3_tri_11;
  reg                 _zz_readLogic_3_tri_12;
  reg                 _zz_readLogic_3_tri_13;
  reg                 _zz_readLogic_3_tri_14;
  reg                 _zz_readLogic_3_tri_15;
  reg                 _zz_readLogic_3_tri_16;
  reg                 _zz_readLogic_3_tri_17;
  reg                 _zz_readLogic_3_tri_18;
  reg                 _zz_readLogic_3_tri_19;
  reg                 _zz_readLogic_3_tri_20;
  reg                 _zz_readLogic_3_tri_21;
  reg                 _zz_readLogic_3_tri_22;
  reg                 _zz_readLogic_3_tri_23;
  reg                 _zz_readLogic_3_tri_24;
  reg                 _zz_readLogic_3_tri_25;
  reg                 _zz_readLogic_3_tri_26;
  reg                 _zz_readLogic_3_tri_27;
  reg                 _zz_readLogic_3_tri_28;
  reg                 _zz_readLogic_3_tri_29;
  reg                 _zz_readLogic_3_tri_30;
  reg                 _zz_readLogic_3_tri_31;
  reg                 _zz_readLogic_3_tri_32;
  reg                 _zz_readLogic_3_tri_33;
  reg                 _zz_readLogic_3_tri_34;
  reg                 _zz_readLogic_3_tri_35;
  reg                 _zz_readLogic_3_tri_36;
  reg                 _zz_readLogic_3_tri_37;
  reg                 _zz_readLogic_3_tri_38;
  reg                 _zz_readLogic_3_tri_39;
  reg                 _zz_readLogic_3_tri_40;
  reg                 _zz_readLogic_3_tri_41;
  reg                 _zz_readLogic_3_tri_42;
  reg                 _zz_readLogic_3_tri_43;
  reg                 _zz_readLogic_3_tri_44;
  reg                 _zz_readLogic_3_tri_45;
  reg                 _zz_readLogic_3_tri_46;
  reg                 _zz_readLogic_3_tri_47;
  reg                 _zz_readLogic_3_tri_48;
  reg                 _zz_readLogic_3_tri_49;
  reg                 _zz_readLogic_3_tri_50;
  reg                 _zz_readLogic_3_tri_51;
  reg                 _zz_readLogic_3_tri_52;
  reg                 _zz_readLogic_3_tri_53;
  reg                 _zz_readLogic_3_tri_54;
  reg                 _zz_readLogic_3_tri_55;
  reg                 _zz_readLogic_3_tri_56;
  reg                 _zz_readLogic_3_tri_57;
  reg                 _zz_readLogic_3_tri_58;
  reg                 _zz_readLogic_3_tri_59;
  reg                 _zz_readLogic_3_tri_60;
  reg                 _zz_readLogic_3_tri_61;
  reg                 _zz_readLogic_3_tri_62;
  reg                 _zz_readLogic_3_tri_63;
  reg                 _zz_readLogic_2_tri;
  reg                 _zz_readLogic_2_tri_1;
  reg                 _zz_readLogic_2_tri_2;
  reg                 _zz_readLogic_2_tri_3;
  reg                 _zz_readLogic_2_tri_4;
  reg                 _zz_readLogic_2_tri_5;
  reg                 _zz_readLogic_2_tri_6;
  reg                 _zz_readLogic_2_tri_7;
  reg                 _zz_readLogic_2_tri_8;
  reg                 _zz_readLogic_2_tri_9;
  reg                 _zz_readLogic_2_tri_10;
  reg                 _zz_readLogic_2_tri_11;
  reg                 _zz_readLogic_2_tri_12;
  reg                 _zz_readLogic_2_tri_13;
  reg                 _zz_readLogic_2_tri_14;
  reg                 _zz_readLogic_2_tri_15;
  reg                 _zz_readLogic_2_tri_16;
  reg                 _zz_readLogic_2_tri_17;
  reg                 _zz_readLogic_2_tri_18;
  reg                 _zz_readLogic_2_tri_19;
  reg                 _zz_readLogic_2_tri_20;
  reg                 _zz_readLogic_2_tri_21;
  reg                 _zz_readLogic_2_tri_22;
  reg                 _zz_readLogic_2_tri_23;
  reg                 _zz_readLogic_2_tri_24;
  reg                 _zz_readLogic_2_tri_25;
  reg                 _zz_readLogic_2_tri_26;
  reg                 _zz_readLogic_2_tri_27;
  reg                 _zz_readLogic_2_tri_28;
  reg                 _zz_readLogic_2_tri_29;
  reg                 _zz_readLogic_2_tri_30;
  reg                 _zz_readLogic_2_tri_31;
  reg                 _zz_readLogic_2_tri_32;
  reg                 _zz_readLogic_2_tri_33;
  reg                 _zz_readLogic_2_tri_34;
  reg                 _zz_readLogic_2_tri_35;
  reg                 _zz_readLogic_2_tri_36;
  reg                 _zz_readLogic_2_tri_37;
  reg                 _zz_readLogic_2_tri_38;
  reg                 _zz_readLogic_2_tri_39;
  reg                 _zz_readLogic_2_tri_40;
  reg                 _zz_readLogic_2_tri_41;
  reg                 _zz_readLogic_2_tri_42;
  reg                 _zz_readLogic_2_tri_43;
  reg                 _zz_readLogic_2_tri_44;
  reg                 _zz_readLogic_2_tri_45;
  reg                 _zz_readLogic_2_tri_46;
  reg                 _zz_readLogic_2_tri_47;
  reg                 _zz_readLogic_2_tri_48;
  reg                 _zz_readLogic_2_tri_49;
  reg                 _zz_readLogic_2_tri_50;
  reg                 _zz_readLogic_2_tri_51;
  reg                 _zz_readLogic_2_tri_52;
  reg                 _zz_readLogic_2_tri_53;
  reg                 _zz_readLogic_2_tri_54;
  reg                 _zz_readLogic_2_tri_55;
  reg                 _zz_readLogic_2_tri_56;
  reg                 _zz_readLogic_2_tri_57;
  reg                 _zz_readLogic_2_tri_58;
  reg                 _zz_readLogic_2_tri_59;
  reg                 _zz_readLogic_2_tri_60;
  reg                 _zz_readLogic_2_tri_61;
  reg                 _zz_readLogic_2_tri_62;
  reg                 _zz_readLogic_2_tri_63;
  reg                 _zz_readLogic_1_tri;
  reg                 _zz_readLogic_1_tri_1;
  reg                 _zz_readLogic_1_tri_2;
  reg                 _zz_readLogic_1_tri_3;
  reg                 _zz_readLogic_1_tri_4;
  reg                 _zz_readLogic_1_tri_5;
  reg                 _zz_readLogic_1_tri_6;
  reg                 _zz_readLogic_1_tri_7;
  reg                 _zz_readLogic_1_tri_8;
  reg                 _zz_readLogic_1_tri_9;
  reg                 _zz_readLogic_1_tri_10;
  reg                 _zz_readLogic_1_tri_11;
  reg                 _zz_readLogic_1_tri_12;
  reg                 _zz_readLogic_1_tri_13;
  reg                 _zz_readLogic_1_tri_14;
  reg                 _zz_readLogic_1_tri_15;
  reg                 _zz_readLogic_1_tri_16;
  reg                 _zz_readLogic_1_tri_17;
  reg                 _zz_readLogic_1_tri_18;
  reg                 _zz_readLogic_1_tri_19;
  reg                 _zz_readLogic_1_tri_20;
  reg                 _zz_readLogic_1_tri_21;
  reg                 _zz_readLogic_1_tri_22;
  reg                 _zz_readLogic_1_tri_23;
  reg                 _zz_readLogic_1_tri_24;
  reg                 _zz_readLogic_1_tri_25;
  reg                 _zz_readLogic_1_tri_26;
  reg                 _zz_readLogic_1_tri_27;
  reg                 _zz_readLogic_1_tri_28;
  reg                 _zz_readLogic_1_tri_29;
  reg                 _zz_readLogic_1_tri_30;
  reg                 _zz_readLogic_1_tri_31;
  reg                 _zz_readLogic_1_tri_32;
  reg                 _zz_readLogic_1_tri_33;
  reg                 _zz_readLogic_1_tri_34;
  reg                 _zz_readLogic_1_tri_35;
  reg                 _zz_readLogic_1_tri_36;
  reg                 _zz_readLogic_1_tri_37;
  reg                 _zz_readLogic_1_tri_38;
  reg                 _zz_readLogic_1_tri_39;
  reg                 _zz_readLogic_1_tri_40;
  reg                 _zz_readLogic_1_tri_41;
  reg                 _zz_readLogic_1_tri_42;
  reg                 _zz_readLogic_1_tri_43;
  reg                 _zz_readLogic_1_tri_44;
  reg                 _zz_readLogic_1_tri_45;
  reg                 _zz_readLogic_1_tri_46;
  reg                 _zz_readLogic_1_tri_47;
  reg                 _zz_readLogic_1_tri_48;
  reg                 _zz_readLogic_1_tri_49;
  reg                 _zz_readLogic_1_tri_50;
  reg                 _zz_readLogic_1_tri_51;
  reg                 _zz_readLogic_1_tri_52;
  reg                 _zz_readLogic_1_tri_53;
  reg                 _zz_readLogic_1_tri_54;
  reg                 _zz_readLogic_1_tri_55;
  reg                 _zz_readLogic_1_tri_56;
  reg                 _zz_readLogic_1_tri_57;
  reg                 _zz_readLogic_1_tri_58;
  reg                 _zz_readLogic_1_tri_59;
  reg                 _zz_readLogic_1_tri_60;
  reg                 _zz_readLogic_1_tri_61;
  reg                 _zz_readLogic_1_tri_62;
  reg                 _zz_readLogic_1_tri_63;
  reg                 _zz_readLogic_0_tri;
  reg                 _zz_readLogic_0_tri_1;
  reg                 _zz_readLogic_0_tri_2;
  reg                 _zz_readLogic_0_tri_3;
  reg                 _zz_readLogic_0_tri_4;
  reg                 _zz_readLogic_0_tri_5;
  reg                 _zz_readLogic_0_tri_6;
  reg                 _zz_readLogic_0_tri_7;
  reg                 _zz_readLogic_0_tri_8;
  reg                 _zz_readLogic_0_tri_9;
  reg                 _zz_readLogic_0_tri_10;
  reg                 _zz_readLogic_0_tri_11;
  reg                 _zz_readLogic_0_tri_12;
  reg                 _zz_readLogic_0_tri_13;
  reg                 _zz_readLogic_0_tri_14;
  reg                 _zz_readLogic_0_tri_15;
  reg                 _zz_readLogic_0_tri_16;
  reg                 _zz_readLogic_0_tri_17;
  reg                 _zz_readLogic_0_tri_18;
  reg                 _zz_readLogic_0_tri_19;
  reg                 _zz_readLogic_0_tri_20;
  reg                 _zz_readLogic_0_tri_21;
  reg                 _zz_readLogic_0_tri_22;
  reg                 _zz_readLogic_0_tri_23;
  reg                 _zz_readLogic_0_tri_24;
  reg                 _zz_readLogic_0_tri_25;
  reg                 _zz_readLogic_0_tri_26;
  reg                 _zz_readLogic_0_tri_27;
  reg                 _zz_readLogic_0_tri_28;
  reg                 _zz_readLogic_0_tri_29;
  reg                 _zz_readLogic_0_tri_30;
  reg                 _zz_readLogic_0_tri_31;
  reg                 _zz_readLogic_0_tri_32;
  reg                 _zz_readLogic_0_tri_33;
  reg                 _zz_readLogic_0_tri_34;
  reg                 _zz_readLogic_0_tri_35;
  reg                 _zz_readLogic_0_tri_36;
  reg                 _zz_readLogic_0_tri_37;
  reg                 _zz_readLogic_0_tri_38;
  reg                 _zz_readLogic_0_tri_39;
  reg                 _zz_readLogic_0_tri_40;
  reg                 _zz_readLogic_0_tri_41;
  reg                 _zz_readLogic_0_tri_42;
  reg                 _zz_readLogic_0_tri_43;
  reg                 _zz_readLogic_0_tri_44;
  reg                 _zz_readLogic_0_tri_45;
  reg                 _zz_readLogic_0_tri_46;
  reg                 _zz_readLogic_0_tri_47;
  reg                 _zz_readLogic_0_tri_48;
  reg                 _zz_readLogic_0_tri_49;
  reg                 _zz_readLogic_0_tri_50;
  reg                 _zz_readLogic_0_tri_51;
  reg                 _zz_readLogic_0_tri_52;
  reg                 _zz_readLogic_0_tri_53;
  reg                 _zz_readLogic_0_tri_54;
  reg                 _zz_readLogic_0_tri_55;
  reg                 _zz_readLogic_0_tri_56;
  reg                 _zz_readLogic_0_tri_57;
  reg                 _zz_readLogic_0_tri_58;
  reg                 _zz_readLogic_0_tri_59;
  reg                 _zz_readLogic_0_tri_60;
  reg                 _zz_readLogic_0_tri_61;
  reg                 _zz_readLogic_0_tri_62;
  reg                 _zz_readLogic_0_tri_63;
  reg        [31:0]   writeFrontend_buffers_0;
  reg        [31:0]   writeFrontend_buffers_1;
  wire       [1:0]    latches_0_write_mask;
  reg        [1:0]    latches_0_write_maskReg;
  reg                 latches_0_write_validReg;
  wire       [31:0]   latches_0_write_data;
  wire                latches_0_write_sample;
  reg        [31:0]   latches_0_storage;
  wire       [1:0]    latches_1_write_mask;
  reg        [1:0]    latches_1_write_maskReg;
  reg                 latches_1_write_validReg;
  wire       [31:0]   latches_1_write_data;
  wire                latches_1_write_sample;
  reg        [31:0]   latches_1_storage;
  wire       [1:0]    latches_2_write_mask;
  reg        [1:0]    latches_2_write_maskReg;
  reg                 latches_2_write_validReg;
  wire       [31:0]   latches_2_write_data;
  wire                latches_2_write_sample;
  reg        [31:0]   latches_2_storage;
  wire       [1:0]    latches_3_write_mask;
  reg        [1:0]    latches_3_write_maskReg;
  reg                 latches_3_write_validReg;
  wire       [31:0]   latches_3_write_data;
  wire                latches_3_write_sample;
  reg        [31:0]   latches_3_storage;
  wire       [1:0]    latches_4_write_mask;
  reg        [1:0]    latches_4_write_maskReg;
  reg                 latches_4_write_validReg;
  wire       [31:0]   latches_4_write_data;
  wire                latches_4_write_sample;
  reg        [31:0]   latches_4_storage;
  wire       [1:0]    latches_5_write_mask;
  reg        [1:0]    latches_5_write_maskReg;
  reg                 latches_5_write_validReg;
  wire       [31:0]   latches_5_write_data;
  wire                latches_5_write_sample;
  reg        [31:0]   latches_5_storage;
  wire       [1:0]    latches_6_write_mask;
  reg        [1:0]    latches_6_write_maskReg;
  reg                 latches_6_write_validReg;
  wire       [31:0]   latches_6_write_data;
  wire                latches_6_write_sample;
  reg        [31:0]   latches_6_storage;
  wire       [1:0]    latches_7_write_mask;
  reg        [1:0]    latches_7_write_maskReg;
  reg                 latches_7_write_validReg;
  wire       [31:0]   latches_7_write_data;
  wire                latches_7_write_sample;
  reg        [31:0]   latches_7_storage;
  wire       [1:0]    latches_8_write_mask;
  reg        [1:0]    latches_8_write_maskReg;
  reg                 latches_8_write_validReg;
  wire       [31:0]   latches_8_write_data;
  wire                latches_8_write_sample;
  reg        [31:0]   latches_8_storage;
  wire       [1:0]    latches_9_write_mask;
  reg        [1:0]    latches_9_write_maskReg;
  reg                 latches_9_write_validReg;
  wire       [31:0]   latches_9_write_data;
  wire                latches_9_write_sample;
  reg        [31:0]   latches_9_storage;
  wire       [1:0]    latches_10_write_mask;
  reg        [1:0]    latches_10_write_maskReg;
  reg                 latches_10_write_validReg;
  wire       [31:0]   latches_10_write_data;
  wire                latches_10_write_sample;
  reg        [31:0]   latches_10_storage;
  wire       [1:0]    latches_11_write_mask;
  reg        [1:0]    latches_11_write_maskReg;
  reg                 latches_11_write_validReg;
  wire       [31:0]   latches_11_write_data;
  wire                latches_11_write_sample;
  reg        [31:0]   latches_11_storage;
  wire       [1:0]    latches_12_write_mask;
  reg        [1:0]    latches_12_write_maskReg;
  reg                 latches_12_write_validReg;
  wire       [31:0]   latches_12_write_data;
  wire                latches_12_write_sample;
  reg        [31:0]   latches_12_storage;
  wire       [1:0]    latches_13_write_mask;
  reg        [1:0]    latches_13_write_maskReg;
  reg                 latches_13_write_validReg;
  wire       [31:0]   latches_13_write_data;
  wire                latches_13_write_sample;
  reg        [31:0]   latches_13_storage;
  wire       [1:0]    latches_14_write_mask;
  reg        [1:0]    latches_14_write_maskReg;
  reg                 latches_14_write_validReg;
  wire       [31:0]   latches_14_write_data;
  wire                latches_14_write_sample;
  reg        [31:0]   latches_14_storage;
  wire       [1:0]    latches_15_write_mask;
  reg        [1:0]    latches_15_write_maskReg;
  reg                 latches_15_write_validReg;
  wire       [31:0]   latches_15_write_data;
  wire                latches_15_write_sample;
  reg        [31:0]   latches_15_storage;
  wire       [1:0]    latches_16_write_mask;
  reg        [1:0]    latches_16_write_maskReg;
  reg                 latches_16_write_validReg;
  wire       [31:0]   latches_16_write_data;
  wire                latches_16_write_sample;
  reg        [31:0]   latches_16_storage;
  wire       [1:0]    latches_17_write_mask;
  reg        [1:0]    latches_17_write_maskReg;
  reg                 latches_17_write_validReg;
  wire       [31:0]   latches_17_write_data;
  wire                latches_17_write_sample;
  reg        [31:0]   latches_17_storage;
  wire       [1:0]    latches_18_write_mask;
  reg        [1:0]    latches_18_write_maskReg;
  reg                 latches_18_write_validReg;
  wire       [31:0]   latches_18_write_data;
  wire                latches_18_write_sample;
  reg        [31:0]   latches_18_storage;
  wire       [1:0]    latches_19_write_mask;
  reg        [1:0]    latches_19_write_maskReg;
  reg                 latches_19_write_validReg;
  wire       [31:0]   latches_19_write_data;
  wire                latches_19_write_sample;
  reg        [31:0]   latches_19_storage;
  wire       [1:0]    latches_20_write_mask;
  reg        [1:0]    latches_20_write_maskReg;
  reg                 latches_20_write_validReg;
  wire       [31:0]   latches_20_write_data;
  wire                latches_20_write_sample;
  reg        [31:0]   latches_20_storage;
  wire       [1:0]    latches_21_write_mask;
  reg        [1:0]    latches_21_write_maskReg;
  reg                 latches_21_write_validReg;
  wire       [31:0]   latches_21_write_data;
  wire                latches_21_write_sample;
  reg        [31:0]   latches_21_storage;
  wire       [1:0]    latches_22_write_mask;
  reg        [1:0]    latches_22_write_maskReg;
  reg                 latches_22_write_validReg;
  wire       [31:0]   latches_22_write_data;
  wire                latches_22_write_sample;
  reg        [31:0]   latches_22_storage;
  wire       [1:0]    latches_23_write_mask;
  reg        [1:0]    latches_23_write_maskReg;
  reg                 latches_23_write_validReg;
  wire       [31:0]   latches_23_write_data;
  wire                latches_23_write_sample;
  reg        [31:0]   latches_23_storage;
  wire       [1:0]    latches_24_write_mask;
  reg        [1:0]    latches_24_write_maskReg;
  reg                 latches_24_write_validReg;
  wire       [31:0]   latches_24_write_data;
  wire                latches_24_write_sample;
  reg        [31:0]   latches_24_storage;
  wire       [1:0]    latches_25_write_mask;
  reg        [1:0]    latches_25_write_maskReg;
  reg                 latches_25_write_validReg;
  wire       [31:0]   latches_25_write_data;
  wire                latches_25_write_sample;
  reg        [31:0]   latches_25_storage;
  wire       [1:0]    latches_26_write_mask;
  reg        [1:0]    latches_26_write_maskReg;
  reg                 latches_26_write_validReg;
  wire       [31:0]   latches_26_write_data;
  wire                latches_26_write_sample;
  reg        [31:0]   latches_26_storage;
  wire       [1:0]    latches_27_write_mask;
  reg        [1:0]    latches_27_write_maskReg;
  reg                 latches_27_write_validReg;
  wire       [31:0]   latches_27_write_data;
  wire                latches_27_write_sample;
  reg        [31:0]   latches_27_storage;
  wire       [1:0]    latches_28_write_mask;
  reg        [1:0]    latches_28_write_maskReg;
  reg                 latches_28_write_validReg;
  wire       [31:0]   latches_28_write_data;
  wire                latches_28_write_sample;
  reg        [31:0]   latches_28_storage;
  wire       [1:0]    latches_29_write_mask;
  reg        [1:0]    latches_29_write_maskReg;
  reg                 latches_29_write_validReg;
  wire       [31:0]   latches_29_write_data;
  wire                latches_29_write_sample;
  reg        [31:0]   latches_29_storage;
  wire       [1:0]    latches_30_write_mask;
  reg        [1:0]    latches_30_write_maskReg;
  reg                 latches_30_write_validReg;
  wire       [31:0]   latches_30_write_data;
  wire                latches_30_write_sample;
  reg        [31:0]   latches_30_storage;
  wire       [1:0]    latches_31_write_mask;
  reg        [1:0]    latches_31_write_maskReg;
  reg                 latches_31_write_validReg;
  wire       [31:0]   latches_31_write_data;
  wire                latches_31_write_sample;
  reg        [31:0]   latches_31_storage;
  wire       [1:0]    latches_32_write_mask;
  reg        [1:0]    latches_32_write_maskReg;
  reg                 latches_32_write_validReg;
  wire       [31:0]   latches_32_write_data;
  wire                latches_32_write_sample;
  reg        [31:0]   latches_32_storage;
  wire       [1:0]    latches_33_write_mask;
  reg        [1:0]    latches_33_write_maskReg;
  reg                 latches_33_write_validReg;
  wire       [31:0]   latches_33_write_data;
  wire                latches_33_write_sample;
  reg        [31:0]   latches_33_storage;
  wire       [1:0]    latches_34_write_mask;
  reg        [1:0]    latches_34_write_maskReg;
  reg                 latches_34_write_validReg;
  wire       [31:0]   latches_34_write_data;
  wire                latches_34_write_sample;
  reg        [31:0]   latches_34_storage;
  wire       [1:0]    latches_35_write_mask;
  reg        [1:0]    latches_35_write_maskReg;
  reg                 latches_35_write_validReg;
  wire       [31:0]   latches_35_write_data;
  wire                latches_35_write_sample;
  reg        [31:0]   latches_35_storage;
  wire       [1:0]    latches_36_write_mask;
  reg        [1:0]    latches_36_write_maskReg;
  reg                 latches_36_write_validReg;
  wire       [31:0]   latches_36_write_data;
  wire                latches_36_write_sample;
  reg        [31:0]   latches_36_storage;
  wire       [1:0]    latches_37_write_mask;
  reg        [1:0]    latches_37_write_maskReg;
  reg                 latches_37_write_validReg;
  wire       [31:0]   latches_37_write_data;
  wire                latches_37_write_sample;
  reg        [31:0]   latches_37_storage;
  wire       [1:0]    latches_38_write_mask;
  reg        [1:0]    latches_38_write_maskReg;
  reg                 latches_38_write_validReg;
  wire       [31:0]   latches_38_write_data;
  wire                latches_38_write_sample;
  reg        [31:0]   latches_38_storage;
  wire       [1:0]    latches_39_write_mask;
  reg        [1:0]    latches_39_write_maskReg;
  reg                 latches_39_write_validReg;
  wire       [31:0]   latches_39_write_data;
  wire                latches_39_write_sample;
  reg        [31:0]   latches_39_storage;
  wire       [1:0]    latches_40_write_mask;
  reg        [1:0]    latches_40_write_maskReg;
  reg                 latches_40_write_validReg;
  wire       [31:0]   latches_40_write_data;
  wire                latches_40_write_sample;
  reg        [31:0]   latches_40_storage;
  wire       [1:0]    latches_41_write_mask;
  reg        [1:0]    latches_41_write_maskReg;
  reg                 latches_41_write_validReg;
  wire       [31:0]   latches_41_write_data;
  wire                latches_41_write_sample;
  reg        [31:0]   latches_41_storage;
  wire       [1:0]    latches_42_write_mask;
  reg        [1:0]    latches_42_write_maskReg;
  reg                 latches_42_write_validReg;
  wire       [31:0]   latches_42_write_data;
  wire                latches_42_write_sample;
  reg        [31:0]   latches_42_storage;
  wire       [1:0]    latches_43_write_mask;
  reg        [1:0]    latches_43_write_maskReg;
  reg                 latches_43_write_validReg;
  wire       [31:0]   latches_43_write_data;
  wire                latches_43_write_sample;
  reg        [31:0]   latches_43_storage;
  wire       [1:0]    latches_44_write_mask;
  reg        [1:0]    latches_44_write_maskReg;
  reg                 latches_44_write_validReg;
  wire       [31:0]   latches_44_write_data;
  wire                latches_44_write_sample;
  reg        [31:0]   latches_44_storage;
  wire       [1:0]    latches_45_write_mask;
  reg        [1:0]    latches_45_write_maskReg;
  reg                 latches_45_write_validReg;
  wire       [31:0]   latches_45_write_data;
  wire                latches_45_write_sample;
  reg        [31:0]   latches_45_storage;
  wire       [1:0]    latches_46_write_mask;
  reg        [1:0]    latches_46_write_maskReg;
  reg                 latches_46_write_validReg;
  wire       [31:0]   latches_46_write_data;
  wire                latches_46_write_sample;
  reg        [31:0]   latches_46_storage;
  wire       [1:0]    latches_47_write_mask;
  reg        [1:0]    latches_47_write_maskReg;
  reg                 latches_47_write_validReg;
  wire       [31:0]   latches_47_write_data;
  wire                latches_47_write_sample;
  reg        [31:0]   latches_47_storage;
  wire       [1:0]    latches_48_write_mask;
  reg        [1:0]    latches_48_write_maskReg;
  reg                 latches_48_write_validReg;
  wire       [31:0]   latches_48_write_data;
  wire                latches_48_write_sample;
  reg        [31:0]   latches_48_storage;
  wire       [1:0]    latches_49_write_mask;
  reg        [1:0]    latches_49_write_maskReg;
  reg                 latches_49_write_validReg;
  wire       [31:0]   latches_49_write_data;
  wire                latches_49_write_sample;
  reg        [31:0]   latches_49_storage;
  wire       [1:0]    latches_50_write_mask;
  reg        [1:0]    latches_50_write_maskReg;
  reg                 latches_50_write_validReg;
  wire       [31:0]   latches_50_write_data;
  wire                latches_50_write_sample;
  reg        [31:0]   latches_50_storage;
  wire       [1:0]    latches_51_write_mask;
  reg        [1:0]    latches_51_write_maskReg;
  reg                 latches_51_write_validReg;
  wire       [31:0]   latches_51_write_data;
  wire                latches_51_write_sample;
  reg        [31:0]   latches_51_storage;
  wire       [1:0]    latches_52_write_mask;
  reg        [1:0]    latches_52_write_maskReg;
  reg                 latches_52_write_validReg;
  wire       [31:0]   latches_52_write_data;
  wire                latches_52_write_sample;
  reg        [31:0]   latches_52_storage;
  wire       [1:0]    latches_53_write_mask;
  reg        [1:0]    latches_53_write_maskReg;
  reg                 latches_53_write_validReg;
  wire       [31:0]   latches_53_write_data;
  wire                latches_53_write_sample;
  reg        [31:0]   latches_53_storage;
  wire       [1:0]    latches_54_write_mask;
  reg        [1:0]    latches_54_write_maskReg;
  reg                 latches_54_write_validReg;
  wire       [31:0]   latches_54_write_data;
  wire                latches_54_write_sample;
  reg        [31:0]   latches_54_storage;
  wire       [1:0]    latches_55_write_mask;
  reg        [1:0]    latches_55_write_maskReg;
  reg                 latches_55_write_validReg;
  wire       [31:0]   latches_55_write_data;
  wire                latches_55_write_sample;
  reg        [31:0]   latches_55_storage;
  wire       [1:0]    latches_56_write_mask;
  reg        [1:0]    latches_56_write_maskReg;
  reg                 latches_56_write_validReg;
  wire       [31:0]   latches_56_write_data;
  wire                latches_56_write_sample;
  reg        [31:0]   latches_56_storage;
  wire       [1:0]    latches_57_write_mask;
  reg        [1:0]    latches_57_write_maskReg;
  reg                 latches_57_write_validReg;
  wire       [31:0]   latches_57_write_data;
  wire                latches_57_write_sample;
  reg        [31:0]   latches_57_storage;
  wire       [1:0]    latches_58_write_mask;
  reg        [1:0]    latches_58_write_maskReg;
  reg                 latches_58_write_validReg;
  wire       [31:0]   latches_58_write_data;
  wire                latches_58_write_sample;
  reg        [31:0]   latches_58_storage;
  wire       [1:0]    latches_59_write_mask;
  reg        [1:0]    latches_59_write_maskReg;
  reg                 latches_59_write_validReg;
  wire       [31:0]   latches_59_write_data;
  wire                latches_59_write_sample;
  reg        [31:0]   latches_59_storage;
  wire       [1:0]    latches_60_write_mask;
  reg        [1:0]    latches_60_write_maskReg;
  reg                 latches_60_write_validReg;
  wire       [31:0]   latches_60_write_data;
  wire                latches_60_write_sample;
  reg        [31:0]   latches_60_storage;
  wire       [1:0]    latches_61_write_mask;
  reg        [1:0]    latches_61_write_maskReg;
  reg                 latches_61_write_validReg;
  wire       [31:0]   latches_61_write_data;
  wire                latches_61_write_sample;
  reg        [31:0]   latches_61_storage;
  wire       [1:0]    latches_62_write_mask;
  reg        [1:0]    latches_62_write_maskReg;
  reg                 latches_62_write_validReg;
  wire       [31:0]   latches_62_write_data;
  wire                latches_62_write_sample;
  reg        [31:0]   latches_62_storage;
  wire       [63:0]   readLogic_0_oh;
  wire       [31:0]   readLogic_0_tri;
  wire       [63:0]   _zz_1;
  wire       [63:0]   readLogic_1_oh;
  wire       [31:0]   readLogic_1_tri;
  wire       [63:0]   _zz_2;
  wire       [63:0]   readLogic_2_oh;
  wire       [31:0]   readLogic_2_tri;
  wire       [63:0]   _zz_3;
  wire       [63:0]   readLogic_3_oh;
  wire       [31:0]   readLogic_3_tri;
  wire       [63:0]   _zz_4;

  assign _zz_readLogic_0_tri_64 = 32'h00000000;
  assign _zz_readLogic_1_tri_64 = 32'h00000000;
  assign _zz_readLogic_2_tri_64 = 32'h00000000;
  assign _zz_readLogic_3_tri_64 = 32'h00000000;
  assign readLogic_0_tri = _zz_readLogic_0_tri_63 ? _zz_readLogic_0_tri_64[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_62 ? latches_0_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_61 ? latches_1_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_60 ? latches_2_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_59 ? latches_3_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_58 ? latches_4_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_57 ? latches_5_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_56 ? latches_6_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_55 ? latches_7_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_54 ? latches_8_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_53 ? latches_9_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_52 ? latches_10_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_51 ? latches_11_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_50 ? latches_12_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_49 ? latches_13_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_48 ? latches_14_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_47 ? latches_15_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_46 ? latches_16_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_45 ? latches_17_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_44 ? latches_18_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_43 ? latches_19_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_42 ? latches_20_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_41 ? latches_21_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_40 ? latches_22_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_39 ? latches_23_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_38 ? latches_24_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_37 ? latches_25_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_36 ? latches_26_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_35 ? latches_27_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_34 ? latches_28_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_33 ? latches_29_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_32 ? latches_30_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_31 ? latches_31_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_30 ? latches_32_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_29 ? latches_33_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_28 ? latches_34_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_27 ? latches_35_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_26 ? latches_36_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_25 ? latches_37_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_24 ? latches_38_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_23 ? latches_39_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_22 ? latches_40_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_21 ? latches_41_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_20 ? latches_42_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_19 ? latches_43_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_18 ? latches_44_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_17 ? latches_45_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_16 ? latches_46_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_15 ? latches_47_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_14 ? latches_48_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_13 ? latches_49_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_12 ? latches_50_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_11 ? latches_51_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_10 ? latches_52_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_9 ? latches_53_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_8 ? latches_54_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_7 ? latches_55_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_6 ? latches_56_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_5 ? latches_57_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_4 ? latches_58_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_3 ? latches_59_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_2 ? latches_60_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri_1 ? latches_61_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_0_tri = _zz_readLogic_0_tri ? latches_62_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_63 ? _zz_readLogic_1_tri_64[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_62 ? latches_0_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_61 ? latches_1_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_60 ? latches_2_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_59 ? latches_3_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_58 ? latches_4_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_57 ? latches_5_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_56 ? latches_6_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_55 ? latches_7_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_54 ? latches_8_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_53 ? latches_9_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_52 ? latches_10_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_51 ? latches_11_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_50 ? latches_12_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_49 ? latches_13_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_48 ? latches_14_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_47 ? latches_15_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_46 ? latches_16_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_45 ? latches_17_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_44 ? latches_18_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_43 ? latches_19_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_42 ? latches_20_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_41 ? latches_21_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_40 ? latches_22_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_39 ? latches_23_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_38 ? latches_24_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_37 ? latches_25_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_36 ? latches_26_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_35 ? latches_27_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_34 ? latches_28_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_33 ? latches_29_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_32 ? latches_30_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_31 ? latches_31_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_30 ? latches_32_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_29 ? latches_33_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_28 ? latches_34_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_27 ? latches_35_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_26 ? latches_36_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_25 ? latches_37_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_24 ? latches_38_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_23 ? latches_39_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_22 ? latches_40_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_21 ? latches_41_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_20 ? latches_42_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_19 ? latches_43_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_18 ? latches_44_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_17 ? latches_45_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_16 ? latches_46_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_15 ? latches_47_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_14 ? latches_48_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_13 ? latches_49_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_12 ? latches_50_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_11 ? latches_51_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_10 ? latches_52_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_9 ? latches_53_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_8 ? latches_54_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_7 ? latches_55_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_6 ? latches_56_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_5 ? latches_57_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_4 ? latches_58_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_3 ? latches_59_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_2 ? latches_60_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri_1 ? latches_61_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_1_tri = _zz_readLogic_1_tri ? latches_62_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_63 ? _zz_readLogic_2_tri_64[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_62 ? latches_0_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_61 ? latches_1_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_60 ? latches_2_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_59 ? latches_3_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_58 ? latches_4_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_57 ? latches_5_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_56 ? latches_6_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_55 ? latches_7_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_54 ? latches_8_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_53 ? latches_9_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_52 ? latches_10_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_51 ? latches_11_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_50 ? latches_12_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_49 ? latches_13_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_48 ? latches_14_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_47 ? latches_15_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_46 ? latches_16_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_45 ? latches_17_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_44 ? latches_18_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_43 ? latches_19_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_42 ? latches_20_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_41 ? latches_21_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_40 ? latches_22_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_39 ? latches_23_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_38 ? latches_24_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_37 ? latches_25_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_36 ? latches_26_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_35 ? latches_27_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_34 ? latches_28_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_33 ? latches_29_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_32 ? latches_30_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_31 ? latches_31_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_30 ? latches_32_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_29 ? latches_33_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_28 ? latches_34_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_27 ? latches_35_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_26 ? latches_36_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_25 ? latches_37_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_24 ? latches_38_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_23 ? latches_39_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_22 ? latches_40_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_21 ? latches_41_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_20 ? latches_42_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_19 ? latches_43_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_18 ? latches_44_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_17 ? latches_45_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_16 ? latches_46_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_15 ? latches_47_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_14 ? latches_48_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_13 ? latches_49_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_12 ? latches_50_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_11 ? latches_51_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_10 ? latches_52_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_9 ? latches_53_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_8 ? latches_54_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_7 ? latches_55_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_6 ? latches_56_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_5 ? latches_57_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_4 ? latches_58_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_3 ? latches_59_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_2 ? latches_60_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri_1 ? latches_61_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_2_tri = _zz_readLogic_2_tri ? latches_62_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_63 ? _zz_readLogic_3_tri_64[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_62 ? latches_0_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_61 ? latches_1_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_60 ? latches_2_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_59 ? latches_3_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_58 ? latches_4_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_57 ? latches_5_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_56 ? latches_6_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_55 ? latches_7_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_54 ? latches_8_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_53 ? latches_9_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_52 ? latches_10_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_51 ? latches_11_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_50 ? latches_12_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_49 ? latches_13_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_48 ? latches_14_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_47 ? latches_15_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_46 ? latches_16_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_45 ? latches_17_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_44 ? latches_18_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_43 ? latches_19_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_42 ? latches_20_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_41 ? latches_21_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_40 ? latches_22_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_39 ? latches_23_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_38 ? latches_24_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_37 ? latches_25_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_36 ? latches_26_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_35 ? latches_27_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_34 ? latches_28_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_33 ? latches_29_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_32 ? latches_30_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_31 ? latches_31_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_30 ? latches_32_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_29 ? latches_33_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_28 ? latches_34_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_27 ? latches_35_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_26 ? latches_36_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_25 ? latches_37_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_24 ? latches_38_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_23 ? latches_39_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_22 ? latches_40_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_21 ? latches_41_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_20 ? latches_42_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_19 ? latches_43_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_18 ? latches_44_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_17 ? latches_45_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_16 ? latches_46_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_15 ? latches_47_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_14 ? latches_48_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_13 ? latches_49_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_12 ? latches_50_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_11 ? latches_51_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_10 ? latches_52_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_9 ? latches_53_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_8 ? latches_54_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_7 ? latches_55_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_6 ? latches_56_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_5 ? latches_57_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_4 ? latches_58_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_3 ? latches_59_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_2 ? latches_60_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri_1 ? latches_61_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  assign readLogic_3_tri = _zz_readLogic_3_tri ? latches_62_storage[31 : 0] : 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
  always @(*) begin
    _zz_readLogic_3_tri = 1'b0;
    if(_zz_4[63]) begin
      _zz_readLogic_3_tri = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_1 = 1'b0;
    if(_zz_4[62]) begin
      _zz_readLogic_3_tri_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_2 = 1'b0;
    if(_zz_4[61]) begin
      _zz_readLogic_3_tri_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_3 = 1'b0;
    if(_zz_4[60]) begin
      _zz_readLogic_3_tri_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_4 = 1'b0;
    if(_zz_4[59]) begin
      _zz_readLogic_3_tri_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_5 = 1'b0;
    if(_zz_4[58]) begin
      _zz_readLogic_3_tri_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_6 = 1'b0;
    if(_zz_4[57]) begin
      _zz_readLogic_3_tri_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_7 = 1'b0;
    if(_zz_4[56]) begin
      _zz_readLogic_3_tri_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_8 = 1'b0;
    if(_zz_4[55]) begin
      _zz_readLogic_3_tri_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_9 = 1'b0;
    if(_zz_4[54]) begin
      _zz_readLogic_3_tri_9 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_10 = 1'b0;
    if(_zz_4[53]) begin
      _zz_readLogic_3_tri_10 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_11 = 1'b0;
    if(_zz_4[52]) begin
      _zz_readLogic_3_tri_11 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_12 = 1'b0;
    if(_zz_4[51]) begin
      _zz_readLogic_3_tri_12 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_13 = 1'b0;
    if(_zz_4[50]) begin
      _zz_readLogic_3_tri_13 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_14 = 1'b0;
    if(_zz_4[49]) begin
      _zz_readLogic_3_tri_14 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_15 = 1'b0;
    if(_zz_4[48]) begin
      _zz_readLogic_3_tri_15 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_16 = 1'b0;
    if(_zz_4[47]) begin
      _zz_readLogic_3_tri_16 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_17 = 1'b0;
    if(_zz_4[46]) begin
      _zz_readLogic_3_tri_17 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_18 = 1'b0;
    if(_zz_4[45]) begin
      _zz_readLogic_3_tri_18 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_19 = 1'b0;
    if(_zz_4[44]) begin
      _zz_readLogic_3_tri_19 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_20 = 1'b0;
    if(_zz_4[43]) begin
      _zz_readLogic_3_tri_20 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_21 = 1'b0;
    if(_zz_4[42]) begin
      _zz_readLogic_3_tri_21 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_22 = 1'b0;
    if(_zz_4[41]) begin
      _zz_readLogic_3_tri_22 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_23 = 1'b0;
    if(_zz_4[40]) begin
      _zz_readLogic_3_tri_23 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_24 = 1'b0;
    if(_zz_4[39]) begin
      _zz_readLogic_3_tri_24 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_25 = 1'b0;
    if(_zz_4[38]) begin
      _zz_readLogic_3_tri_25 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_26 = 1'b0;
    if(_zz_4[37]) begin
      _zz_readLogic_3_tri_26 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_27 = 1'b0;
    if(_zz_4[36]) begin
      _zz_readLogic_3_tri_27 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_28 = 1'b0;
    if(_zz_4[35]) begin
      _zz_readLogic_3_tri_28 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_29 = 1'b0;
    if(_zz_4[34]) begin
      _zz_readLogic_3_tri_29 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_30 = 1'b0;
    if(_zz_4[33]) begin
      _zz_readLogic_3_tri_30 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_31 = 1'b0;
    if(_zz_4[32]) begin
      _zz_readLogic_3_tri_31 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_32 = 1'b0;
    if(_zz_4[31]) begin
      _zz_readLogic_3_tri_32 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_33 = 1'b0;
    if(_zz_4[30]) begin
      _zz_readLogic_3_tri_33 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_34 = 1'b0;
    if(_zz_4[29]) begin
      _zz_readLogic_3_tri_34 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_35 = 1'b0;
    if(_zz_4[28]) begin
      _zz_readLogic_3_tri_35 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_36 = 1'b0;
    if(_zz_4[27]) begin
      _zz_readLogic_3_tri_36 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_37 = 1'b0;
    if(_zz_4[26]) begin
      _zz_readLogic_3_tri_37 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_38 = 1'b0;
    if(_zz_4[25]) begin
      _zz_readLogic_3_tri_38 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_39 = 1'b0;
    if(_zz_4[24]) begin
      _zz_readLogic_3_tri_39 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_40 = 1'b0;
    if(_zz_4[23]) begin
      _zz_readLogic_3_tri_40 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_41 = 1'b0;
    if(_zz_4[22]) begin
      _zz_readLogic_3_tri_41 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_42 = 1'b0;
    if(_zz_4[21]) begin
      _zz_readLogic_3_tri_42 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_43 = 1'b0;
    if(_zz_4[20]) begin
      _zz_readLogic_3_tri_43 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_44 = 1'b0;
    if(_zz_4[19]) begin
      _zz_readLogic_3_tri_44 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_45 = 1'b0;
    if(_zz_4[18]) begin
      _zz_readLogic_3_tri_45 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_46 = 1'b0;
    if(_zz_4[17]) begin
      _zz_readLogic_3_tri_46 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_47 = 1'b0;
    if(_zz_4[16]) begin
      _zz_readLogic_3_tri_47 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_48 = 1'b0;
    if(_zz_4[15]) begin
      _zz_readLogic_3_tri_48 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_49 = 1'b0;
    if(_zz_4[14]) begin
      _zz_readLogic_3_tri_49 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_50 = 1'b0;
    if(_zz_4[13]) begin
      _zz_readLogic_3_tri_50 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_51 = 1'b0;
    if(_zz_4[12]) begin
      _zz_readLogic_3_tri_51 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_52 = 1'b0;
    if(_zz_4[11]) begin
      _zz_readLogic_3_tri_52 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_53 = 1'b0;
    if(_zz_4[10]) begin
      _zz_readLogic_3_tri_53 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_54 = 1'b0;
    if(_zz_4[9]) begin
      _zz_readLogic_3_tri_54 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_55 = 1'b0;
    if(_zz_4[8]) begin
      _zz_readLogic_3_tri_55 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_56 = 1'b0;
    if(_zz_4[7]) begin
      _zz_readLogic_3_tri_56 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_57 = 1'b0;
    if(_zz_4[6]) begin
      _zz_readLogic_3_tri_57 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_58 = 1'b0;
    if(_zz_4[5]) begin
      _zz_readLogic_3_tri_58 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_59 = 1'b0;
    if(_zz_4[4]) begin
      _zz_readLogic_3_tri_59 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_60 = 1'b0;
    if(_zz_4[3]) begin
      _zz_readLogic_3_tri_60 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_61 = 1'b0;
    if(_zz_4[2]) begin
      _zz_readLogic_3_tri_61 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_62 = 1'b0;
    if(_zz_4[1]) begin
      _zz_readLogic_3_tri_62 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_3_tri_63 = 1'b0;
    if(_zz_4[0]) begin
      _zz_readLogic_3_tri_63 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri = 1'b0;
    if(_zz_3[63]) begin
      _zz_readLogic_2_tri = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_1 = 1'b0;
    if(_zz_3[62]) begin
      _zz_readLogic_2_tri_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_2 = 1'b0;
    if(_zz_3[61]) begin
      _zz_readLogic_2_tri_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_3 = 1'b0;
    if(_zz_3[60]) begin
      _zz_readLogic_2_tri_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_4 = 1'b0;
    if(_zz_3[59]) begin
      _zz_readLogic_2_tri_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_5 = 1'b0;
    if(_zz_3[58]) begin
      _zz_readLogic_2_tri_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_6 = 1'b0;
    if(_zz_3[57]) begin
      _zz_readLogic_2_tri_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_7 = 1'b0;
    if(_zz_3[56]) begin
      _zz_readLogic_2_tri_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_8 = 1'b0;
    if(_zz_3[55]) begin
      _zz_readLogic_2_tri_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_9 = 1'b0;
    if(_zz_3[54]) begin
      _zz_readLogic_2_tri_9 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_10 = 1'b0;
    if(_zz_3[53]) begin
      _zz_readLogic_2_tri_10 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_11 = 1'b0;
    if(_zz_3[52]) begin
      _zz_readLogic_2_tri_11 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_12 = 1'b0;
    if(_zz_3[51]) begin
      _zz_readLogic_2_tri_12 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_13 = 1'b0;
    if(_zz_3[50]) begin
      _zz_readLogic_2_tri_13 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_14 = 1'b0;
    if(_zz_3[49]) begin
      _zz_readLogic_2_tri_14 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_15 = 1'b0;
    if(_zz_3[48]) begin
      _zz_readLogic_2_tri_15 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_16 = 1'b0;
    if(_zz_3[47]) begin
      _zz_readLogic_2_tri_16 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_17 = 1'b0;
    if(_zz_3[46]) begin
      _zz_readLogic_2_tri_17 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_18 = 1'b0;
    if(_zz_3[45]) begin
      _zz_readLogic_2_tri_18 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_19 = 1'b0;
    if(_zz_3[44]) begin
      _zz_readLogic_2_tri_19 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_20 = 1'b0;
    if(_zz_3[43]) begin
      _zz_readLogic_2_tri_20 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_21 = 1'b0;
    if(_zz_3[42]) begin
      _zz_readLogic_2_tri_21 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_22 = 1'b0;
    if(_zz_3[41]) begin
      _zz_readLogic_2_tri_22 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_23 = 1'b0;
    if(_zz_3[40]) begin
      _zz_readLogic_2_tri_23 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_24 = 1'b0;
    if(_zz_3[39]) begin
      _zz_readLogic_2_tri_24 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_25 = 1'b0;
    if(_zz_3[38]) begin
      _zz_readLogic_2_tri_25 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_26 = 1'b0;
    if(_zz_3[37]) begin
      _zz_readLogic_2_tri_26 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_27 = 1'b0;
    if(_zz_3[36]) begin
      _zz_readLogic_2_tri_27 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_28 = 1'b0;
    if(_zz_3[35]) begin
      _zz_readLogic_2_tri_28 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_29 = 1'b0;
    if(_zz_3[34]) begin
      _zz_readLogic_2_tri_29 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_30 = 1'b0;
    if(_zz_3[33]) begin
      _zz_readLogic_2_tri_30 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_31 = 1'b0;
    if(_zz_3[32]) begin
      _zz_readLogic_2_tri_31 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_32 = 1'b0;
    if(_zz_3[31]) begin
      _zz_readLogic_2_tri_32 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_33 = 1'b0;
    if(_zz_3[30]) begin
      _zz_readLogic_2_tri_33 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_34 = 1'b0;
    if(_zz_3[29]) begin
      _zz_readLogic_2_tri_34 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_35 = 1'b0;
    if(_zz_3[28]) begin
      _zz_readLogic_2_tri_35 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_36 = 1'b0;
    if(_zz_3[27]) begin
      _zz_readLogic_2_tri_36 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_37 = 1'b0;
    if(_zz_3[26]) begin
      _zz_readLogic_2_tri_37 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_38 = 1'b0;
    if(_zz_3[25]) begin
      _zz_readLogic_2_tri_38 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_39 = 1'b0;
    if(_zz_3[24]) begin
      _zz_readLogic_2_tri_39 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_40 = 1'b0;
    if(_zz_3[23]) begin
      _zz_readLogic_2_tri_40 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_41 = 1'b0;
    if(_zz_3[22]) begin
      _zz_readLogic_2_tri_41 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_42 = 1'b0;
    if(_zz_3[21]) begin
      _zz_readLogic_2_tri_42 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_43 = 1'b0;
    if(_zz_3[20]) begin
      _zz_readLogic_2_tri_43 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_44 = 1'b0;
    if(_zz_3[19]) begin
      _zz_readLogic_2_tri_44 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_45 = 1'b0;
    if(_zz_3[18]) begin
      _zz_readLogic_2_tri_45 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_46 = 1'b0;
    if(_zz_3[17]) begin
      _zz_readLogic_2_tri_46 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_47 = 1'b0;
    if(_zz_3[16]) begin
      _zz_readLogic_2_tri_47 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_48 = 1'b0;
    if(_zz_3[15]) begin
      _zz_readLogic_2_tri_48 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_49 = 1'b0;
    if(_zz_3[14]) begin
      _zz_readLogic_2_tri_49 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_50 = 1'b0;
    if(_zz_3[13]) begin
      _zz_readLogic_2_tri_50 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_51 = 1'b0;
    if(_zz_3[12]) begin
      _zz_readLogic_2_tri_51 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_52 = 1'b0;
    if(_zz_3[11]) begin
      _zz_readLogic_2_tri_52 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_53 = 1'b0;
    if(_zz_3[10]) begin
      _zz_readLogic_2_tri_53 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_54 = 1'b0;
    if(_zz_3[9]) begin
      _zz_readLogic_2_tri_54 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_55 = 1'b0;
    if(_zz_3[8]) begin
      _zz_readLogic_2_tri_55 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_56 = 1'b0;
    if(_zz_3[7]) begin
      _zz_readLogic_2_tri_56 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_57 = 1'b0;
    if(_zz_3[6]) begin
      _zz_readLogic_2_tri_57 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_58 = 1'b0;
    if(_zz_3[5]) begin
      _zz_readLogic_2_tri_58 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_59 = 1'b0;
    if(_zz_3[4]) begin
      _zz_readLogic_2_tri_59 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_60 = 1'b0;
    if(_zz_3[3]) begin
      _zz_readLogic_2_tri_60 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_61 = 1'b0;
    if(_zz_3[2]) begin
      _zz_readLogic_2_tri_61 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_62 = 1'b0;
    if(_zz_3[1]) begin
      _zz_readLogic_2_tri_62 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_2_tri_63 = 1'b0;
    if(_zz_3[0]) begin
      _zz_readLogic_2_tri_63 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri = 1'b0;
    if(_zz_2[63]) begin
      _zz_readLogic_1_tri = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_1 = 1'b0;
    if(_zz_2[62]) begin
      _zz_readLogic_1_tri_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_2 = 1'b0;
    if(_zz_2[61]) begin
      _zz_readLogic_1_tri_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_3 = 1'b0;
    if(_zz_2[60]) begin
      _zz_readLogic_1_tri_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_4 = 1'b0;
    if(_zz_2[59]) begin
      _zz_readLogic_1_tri_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_5 = 1'b0;
    if(_zz_2[58]) begin
      _zz_readLogic_1_tri_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_6 = 1'b0;
    if(_zz_2[57]) begin
      _zz_readLogic_1_tri_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_7 = 1'b0;
    if(_zz_2[56]) begin
      _zz_readLogic_1_tri_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_8 = 1'b0;
    if(_zz_2[55]) begin
      _zz_readLogic_1_tri_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_9 = 1'b0;
    if(_zz_2[54]) begin
      _zz_readLogic_1_tri_9 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_10 = 1'b0;
    if(_zz_2[53]) begin
      _zz_readLogic_1_tri_10 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_11 = 1'b0;
    if(_zz_2[52]) begin
      _zz_readLogic_1_tri_11 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_12 = 1'b0;
    if(_zz_2[51]) begin
      _zz_readLogic_1_tri_12 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_13 = 1'b0;
    if(_zz_2[50]) begin
      _zz_readLogic_1_tri_13 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_14 = 1'b0;
    if(_zz_2[49]) begin
      _zz_readLogic_1_tri_14 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_15 = 1'b0;
    if(_zz_2[48]) begin
      _zz_readLogic_1_tri_15 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_16 = 1'b0;
    if(_zz_2[47]) begin
      _zz_readLogic_1_tri_16 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_17 = 1'b0;
    if(_zz_2[46]) begin
      _zz_readLogic_1_tri_17 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_18 = 1'b0;
    if(_zz_2[45]) begin
      _zz_readLogic_1_tri_18 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_19 = 1'b0;
    if(_zz_2[44]) begin
      _zz_readLogic_1_tri_19 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_20 = 1'b0;
    if(_zz_2[43]) begin
      _zz_readLogic_1_tri_20 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_21 = 1'b0;
    if(_zz_2[42]) begin
      _zz_readLogic_1_tri_21 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_22 = 1'b0;
    if(_zz_2[41]) begin
      _zz_readLogic_1_tri_22 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_23 = 1'b0;
    if(_zz_2[40]) begin
      _zz_readLogic_1_tri_23 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_24 = 1'b0;
    if(_zz_2[39]) begin
      _zz_readLogic_1_tri_24 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_25 = 1'b0;
    if(_zz_2[38]) begin
      _zz_readLogic_1_tri_25 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_26 = 1'b0;
    if(_zz_2[37]) begin
      _zz_readLogic_1_tri_26 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_27 = 1'b0;
    if(_zz_2[36]) begin
      _zz_readLogic_1_tri_27 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_28 = 1'b0;
    if(_zz_2[35]) begin
      _zz_readLogic_1_tri_28 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_29 = 1'b0;
    if(_zz_2[34]) begin
      _zz_readLogic_1_tri_29 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_30 = 1'b0;
    if(_zz_2[33]) begin
      _zz_readLogic_1_tri_30 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_31 = 1'b0;
    if(_zz_2[32]) begin
      _zz_readLogic_1_tri_31 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_32 = 1'b0;
    if(_zz_2[31]) begin
      _zz_readLogic_1_tri_32 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_33 = 1'b0;
    if(_zz_2[30]) begin
      _zz_readLogic_1_tri_33 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_34 = 1'b0;
    if(_zz_2[29]) begin
      _zz_readLogic_1_tri_34 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_35 = 1'b0;
    if(_zz_2[28]) begin
      _zz_readLogic_1_tri_35 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_36 = 1'b0;
    if(_zz_2[27]) begin
      _zz_readLogic_1_tri_36 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_37 = 1'b0;
    if(_zz_2[26]) begin
      _zz_readLogic_1_tri_37 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_38 = 1'b0;
    if(_zz_2[25]) begin
      _zz_readLogic_1_tri_38 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_39 = 1'b0;
    if(_zz_2[24]) begin
      _zz_readLogic_1_tri_39 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_40 = 1'b0;
    if(_zz_2[23]) begin
      _zz_readLogic_1_tri_40 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_41 = 1'b0;
    if(_zz_2[22]) begin
      _zz_readLogic_1_tri_41 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_42 = 1'b0;
    if(_zz_2[21]) begin
      _zz_readLogic_1_tri_42 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_43 = 1'b0;
    if(_zz_2[20]) begin
      _zz_readLogic_1_tri_43 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_44 = 1'b0;
    if(_zz_2[19]) begin
      _zz_readLogic_1_tri_44 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_45 = 1'b0;
    if(_zz_2[18]) begin
      _zz_readLogic_1_tri_45 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_46 = 1'b0;
    if(_zz_2[17]) begin
      _zz_readLogic_1_tri_46 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_47 = 1'b0;
    if(_zz_2[16]) begin
      _zz_readLogic_1_tri_47 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_48 = 1'b0;
    if(_zz_2[15]) begin
      _zz_readLogic_1_tri_48 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_49 = 1'b0;
    if(_zz_2[14]) begin
      _zz_readLogic_1_tri_49 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_50 = 1'b0;
    if(_zz_2[13]) begin
      _zz_readLogic_1_tri_50 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_51 = 1'b0;
    if(_zz_2[12]) begin
      _zz_readLogic_1_tri_51 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_52 = 1'b0;
    if(_zz_2[11]) begin
      _zz_readLogic_1_tri_52 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_53 = 1'b0;
    if(_zz_2[10]) begin
      _zz_readLogic_1_tri_53 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_54 = 1'b0;
    if(_zz_2[9]) begin
      _zz_readLogic_1_tri_54 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_55 = 1'b0;
    if(_zz_2[8]) begin
      _zz_readLogic_1_tri_55 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_56 = 1'b0;
    if(_zz_2[7]) begin
      _zz_readLogic_1_tri_56 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_57 = 1'b0;
    if(_zz_2[6]) begin
      _zz_readLogic_1_tri_57 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_58 = 1'b0;
    if(_zz_2[5]) begin
      _zz_readLogic_1_tri_58 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_59 = 1'b0;
    if(_zz_2[4]) begin
      _zz_readLogic_1_tri_59 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_60 = 1'b0;
    if(_zz_2[3]) begin
      _zz_readLogic_1_tri_60 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_61 = 1'b0;
    if(_zz_2[2]) begin
      _zz_readLogic_1_tri_61 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_62 = 1'b0;
    if(_zz_2[1]) begin
      _zz_readLogic_1_tri_62 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_1_tri_63 = 1'b0;
    if(_zz_2[0]) begin
      _zz_readLogic_1_tri_63 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri = 1'b0;
    if(_zz_1[63]) begin
      _zz_readLogic_0_tri = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_1 = 1'b0;
    if(_zz_1[62]) begin
      _zz_readLogic_0_tri_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_2 = 1'b0;
    if(_zz_1[61]) begin
      _zz_readLogic_0_tri_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_3 = 1'b0;
    if(_zz_1[60]) begin
      _zz_readLogic_0_tri_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_4 = 1'b0;
    if(_zz_1[59]) begin
      _zz_readLogic_0_tri_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_5 = 1'b0;
    if(_zz_1[58]) begin
      _zz_readLogic_0_tri_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_6 = 1'b0;
    if(_zz_1[57]) begin
      _zz_readLogic_0_tri_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_7 = 1'b0;
    if(_zz_1[56]) begin
      _zz_readLogic_0_tri_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_8 = 1'b0;
    if(_zz_1[55]) begin
      _zz_readLogic_0_tri_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_9 = 1'b0;
    if(_zz_1[54]) begin
      _zz_readLogic_0_tri_9 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_10 = 1'b0;
    if(_zz_1[53]) begin
      _zz_readLogic_0_tri_10 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_11 = 1'b0;
    if(_zz_1[52]) begin
      _zz_readLogic_0_tri_11 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_12 = 1'b0;
    if(_zz_1[51]) begin
      _zz_readLogic_0_tri_12 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_13 = 1'b0;
    if(_zz_1[50]) begin
      _zz_readLogic_0_tri_13 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_14 = 1'b0;
    if(_zz_1[49]) begin
      _zz_readLogic_0_tri_14 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_15 = 1'b0;
    if(_zz_1[48]) begin
      _zz_readLogic_0_tri_15 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_16 = 1'b0;
    if(_zz_1[47]) begin
      _zz_readLogic_0_tri_16 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_17 = 1'b0;
    if(_zz_1[46]) begin
      _zz_readLogic_0_tri_17 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_18 = 1'b0;
    if(_zz_1[45]) begin
      _zz_readLogic_0_tri_18 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_19 = 1'b0;
    if(_zz_1[44]) begin
      _zz_readLogic_0_tri_19 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_20 = 1'b0;
    if(_zz_1[43]) begin
      _zz_readLogic_0_tri_20 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_21 = 1'b0;
    if(_zz_1[42]) begin
      _zz_readLogic_0_tri_21 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_22 = 1'b0;
    if(_zz_1[41]) begin
      _zz_readLogic_0_tri_22 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_23 = 1'b0;
    if(_zz_1[40]) begin
      _zz_readLogic_0_tri_23 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_24 = 1'b0;
    if(_zz_1[39]) begin
      _zz_readLogic_0_tri_24 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_25 = 1'b0;
    if(_zz_1[38]) begin
      _zz_readLogic_0_tri_25 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_26 = 1'b0;
    if(_zz_1[37]) begin
      _zz_readLogic_0_tri_26 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_27 = 1'b0;
    if(_zz_1[36]) begin
      _zz_readLogic_0_tri_27 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_28 = 1'b0;
    if(_zz_1[35]) begin
      _zz_readLogic_0_tri_28 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_29 = 1'b0;
    if(_zz_1[34]) begin
      _zz_readLogic_0_tri_29 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_30 = 1'b0;
    if(_zz_1[33]) begin
      _zz_readLogic_0_tri_30 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_31 = 1'b0;
    if(_zz_1[32]) begin
      _zz_readLogic_0_tri_31 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_32 = 1'b0;
    if(_zz_1[31]) begin
      _zz_readLogic_0_tri_32 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_33 = 1'b0;
    if(_zz_1[30]) begin
      _zz_readLogic_0_tri_33 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_34 = 1'b0;
    if(_zz_1[29]) begin
      _zz_readLogic_0_tri_34 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_35 = 1'b0;
    if(_zz_1[28]) begin
      _zz_readLogic_0_tri_35 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_36 = 1'b0;
    if(_zz_1[27]) begin
      _zz_readLogic_0_tri_36 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_37 = 1'b0;
    if(_zz_1[26]) begin
      _zz_readLogic_0_tri_37 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_38 = 1'b0;
    if(_zz_1[25]) begin
      _zz_readLogic_0_tri_38 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_39 = 1'b0;
    if(_zz_1[24]) begin
      _zz_readLogic_0_tri_39 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_40 = 1'b0;
    if(_zz_1[23]) begin
      _zz_readLogic_0_tri_40 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_41 = 1'b0;
    if(_zz_1[22]) begin
      _zz_readLogic_0_tri_41 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_42 = 1'b0;
    if(_zz_1[21]) begin
      _zz_readLogic_0_tri_42 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_43 = 1'b0;
    if(_zz_1[20]) begin
      _zz_readLogic_0_tri_43 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_44 = 1'b0;
    if(_zz_1[19]) begin
      _zz_readLogic_0_tri_44 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_45 = 1'b0;
    if(_zz_1[18]) begin
      _zz_readLogic_0_tri_45 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_46 = 1'b0;
    if(_zz_1[17]) begin
      _zz_readLogic_0_tri_46 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_47 = 1'b0;
    if(_zz_1[16]) begin
      _zz_readLogic_0_tri_47 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_48 = 1'b0;
    if(_zz_1[15]) begin
      _zz_readLogic_0_tri_48 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_49 = 1'b0;
    if(_zz_1[14]) begin
      _zz_readLogic_0_tri_49 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_50 = 1'b0;
    if(_zz_1[13]) begin
      _zz_readLogic_0_tri_50 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_51 = 1'b0;
    if(_zz_1[12]) begin
      _zz_readLogic_0_tri_51 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_52 = 1'b0;
    if(_zz_1[11]) begin
      _zz_readLogic_0_tri_52 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_53 = 1'b0;
    if(_zz_1[10]) begin
      _zz_readLogic_0_tri_53 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_54 = 1'b0;
    if(_zz_1[9]) begin
      _zz_readLogic_0_tri_54 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_55 = 1'b0;
    if(_zz_1[8]) begin
      _zz_readLogic_0_tri_55 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_56 = 1'b0;
    if(_zz_1[7]) begin
      _zz_readLogic_0_tri_56 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_57 = 1'b0;
    if(_zz_1[6]) begin
      _zz_readLogic_0_tri_57 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_58 = 1'b0;
    if(_zz_1[5]) begin
      _zz_readLogic_0_tri_58 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_59 = 1'b0;
    if(_zz_1[4]) begin
      _zz_readLogic_0_tri_59 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_60 = 1'b0;
    if(_zz_1[3]) begin
      _zz_readLogic_0_tri_60 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_61 = 1'b0;
    if(_zz_1[2]) begin
      _zz_readLogic_0_tri_61 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_62 = 1'b0;
    if(_zz_1[1]) begin
      _zz_readLogic_0_tri_62 = 1'b1;
    end
  end

  always @(*) begin
    _zz_readLogic_0_tri_63 = 1'b0;
    if(_zz_1[0]) begin
      _zz_readLogic_0_tri_63 = 1'b1;
    end
  end

  assign latches_0_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h01)),(io_writes_0_valid && (io_writes_0_address == 6'h01))};
  assign latches_0_write_data = ((latches_0_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_0_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_0_write_sample = ((! clk) && latches_0_write_validReg);
  always @(*) begin
    if(latches_0_write_sample) begin
      latches_0_storage = latches_0_write_data;
    end
  end

  assign latches_1_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h02)),(io_writes_0_valid && (io_writes_0_address == 6'h02))};
  assign latches_1_write_data = ((latches_1_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_1_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_1_write_sample = ((! clk) && latches_1_write_validReg);
  always @(*) begin
    if(latches_1_write_sample) begin
      latches_1_storage = latches_1_write_data;
    end
  end

  assign latches_2_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h03)),(io_writes_0_valid && (io_writes_0_address == 6'h03))};
  assign latches_2_write_data = ((latches_2_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_2_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_2_write_sample = ((! clk) && latches_2_write_validReg);
  always @(*) begin
    if(latches_2_write_sample) begin
      latches_2_storage = latches_2_write_data;
    end
  end

  assign latches_3_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h04)),(io_writes_0_valid && (io_writes_0_address == 6'h04))};
  assign latches_3_write_data = ((latches_3_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_3_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_3_write_sample = ((! clk) && latches_3_write_validReg);
  always @(*) begin
    if(latches_3_write_sample) begin
      latches_3_storage = latches_3_write_data;
    end
  end

  assign latches_4_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h05)),(io_writes_0_valid && (io_writes_0_address == 6'h05))};
  assign latches_4_write_data = ((latches_4_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_4_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_4_write_sample = ((! clk) && latches_4_write_validReg);
  always @(*) begin
    if(latches_4_write_sample) begin
      latches_4_storage = latches_4_write_data;
    end
  end

  assign latches_5_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h06)),(io_writes_0_valid && (io_writes_0_address == 6'h06))};
  assign latches_5_write_data = ((latches_5_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_5_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_5_write_sample = ((! clk) && latches_5_write_validReg);
  always @(*) begin
    if(latches_5_write_sample) begin
      latches_5_storage = latches_5_write_data;
    end
  end

  assign latches_6_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h07)),(io_writes_0_valid && (io_writes_0_address == 6'h07))};
  assign latches_6_write_data = ((latches_6_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_6_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_6_write_sample = ((! clk) && latches_6_write_validReg);
  always @(*) begin
    if(latches_6_write_sample) begin
      latches_6_storage = latches_6_write_data;
    end
  end

  assign latches_7_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h08)),(io_writes_0_valid && (io_writes_0_address == 6'h08))};
  assign latches_7_write_data = ((latches_7_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_7_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_7_write_sample = ((! clk) && latches_7_write_validReg);
  always @(*) begin
    if(latches_7_write_sample) begin
      latches_7_storage = latches_7_write_data;
    end
  end

  assign latches_8_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h09)),(io_writes_0_valid && (io_writes_0_address == 6'h09))};
  assign latches_8_write_data = ((latches_8_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_8_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_8_write_sample = ((! clk) && latches_8_write_validReg);
  always @(*) begin
    if(latches_8_write_sample) begin
      latches_8_storage = latches_8_write_data;
    end
  end

  assign latches_9_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h0a)),(io_writes_0_valid && (io_writes_0_address == 6'h0a))};
  assign latches_9_write_data = ((latches_9_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_9_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_9_write_sample = ((! clk) && latches_9_write_validReg);
  always @(*) begin
    if(latches_9_write_sample) begin
      latches_9_storage = latches_9_write_data;
    end
  end

  assign latches_10_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h0b)),(io_writes_0_valid && (io_writes_0_address == 6'h0b))};
  assign latches_10_write_data = ((latches_10_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_10_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_10_write_sample = ((! clk) && latches_10_write_validReg);
  always @(*) begin
    if(latches_10_write_sample) begin
      latches_10_storage = latches_10_write_data;
    end
  end

  assign latches_11_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h0c)),(io_writes_0_valid && (io_writes_0_address == 6'h0c))};
  assign latches_11_write_data = ((latches_11_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_11_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_11_write_sample = ((! clk) && latches_11_write_validReg);
  always @(*) begin
    if(latches_11_write_sample) begin
      latches_11_storage = latches_11_write_data;
    end
  end

  assign latches_12_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h0d)),(io_writes_0_valid && (io_writes_0_address == 6'h0d))};
  assign latches_12_write_data = ((latches_12_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_12_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_12_write_sample = ((! clk) && latches_12_write_validReg);
  always @(*) begin
    if(latches_12_write_sample) begin
      latches_12_storage = latches_12_write_data;
    end
  end

  assign latches_13_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h0e)),(io_writes_0_valid && (io_writes_0_address == 6'h0e))};
  assign latches_13_write_data = ((latches_13_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_13_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_13_write_sample = ((! clk) && latches_13_write_validReg);
  always @(*) begin
    if(latches_13_write_sample) begin
      latches_13_storage = latches_13_write_data;
    end
  end

  assign latches_14_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h0f)),(io_writes_0_valid && (io_writes_0_address == 6'h0f))};
  assign latches_14_write_data = ((latches_14_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_14_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_14_write_sample = ((! clk) && latches_14_write_validReg);
  always @(*) begin
    if(latches_14_write_sample) begin
      latches_14_storage = latches_14_write_data;
    end
  end

  assign latches_15_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h10)),(io_writes_0_valid && (io_writes_0_address == 6'h10))};
  assign latches_15_write_data = ((latches_15_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_15_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_15_write_sample = ((! clk) && latches_15_write_validReg);
  always @(*) begin
    if(latches_15_write_sample) begin
      latches_15_storage = latches_15_write_data;
    end
  end

  assign latches_16_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h11)),(io_writes_0_valid && (io_writes_0_address == 6'h11))};
  assign latches_16_write_data = ((latches_16_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_16_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_16_write_sample = ((! clk) && latches_16_write_validReg);
  always @(*) begin
    if(latches_16_write_sample) begin
      latches_16_storage = latches_16_write_data;
    end
  end

  assign latches_17_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h12)),(io_writes_0_valid && (io_writes_0_address == 6'h12))};
  assign latches_17_write_data = ((latches_17_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_17_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_17_write_sample = ((! clk) && latches_17_write_validReg);
  always @(*) begin
    if(latches_17_write_sample) begin
      latches_17_storage = latches_17_write_data;
    end
  end

  assign latches_18_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h13)),(io_writes_0_valid && (io_writes_0_address == 6'h13))};
  assign latches_18_write_data = ((latches_18_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_18_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_18_write_sample = ((! clk) && latches_18_write_validReg);
  always @(*) begin
    if(latches_18_write_sample) begin
      latches_18_storage = latches_18_write_data;
    end
  end

  assign latches_19_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h14)),(io_writes_0_valid && (io_writes_0_address == 6'h14))};
  assign latches_19_write_data = ((latches_19_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_19_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_19_write_sample = ((! clk) && latches_19_write_validReg);
  always @(*) begin
    if(latches_19_write_sample) begin
      latches_19_storage = latches_19_write_data;
    end
  end

  assign latches_20_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h15)),(io_writes_0_valid && (io_writes_0_address == 6'h15))};
  assign latches_20_write_data = ((latches_20_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_20_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_20_write_sample = ((! clk) && latches_20_write_validReg);
  always @(*) begin
    if(latches_20_write_sample) begin
      latches_20_storage = latches_20_write_data;
    end
  end

  assign latches_21_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h16)),(io_writes_0_valid && (io_writes_0_address == 6'h16))};
  assign latches_21_write_data = ((latches_21_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_21_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_21_write_sample = ((! clk) && latches_21_write_validReg);
  always @(*) begin
    if(latches_21_write_sample) begin
      latches_21_storage = latches_21_write_data;
    end
  end

  assign latches_22_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h17)),(io_writes_0_valid && (io_writes_0_address == 6'h17))};
  assign latches_22_write_data = ((latches_22_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_22_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_22_write_sample = ((! clk) && latches_22_write_validReg);
  always @(*) begin
    if(latches_22_write_sample) begin
      latches_22_storage = latches_22_write_data;
    end
  end

  assign latches_23_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h18)),(io_writes_0_valid && (io_writes_0_address == 6'h18))};
  assign latches_23_write_data = ((latches_23_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_23_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_23_write_sample = ((! clk) && latches_23_write_validReg);
  always @(*) begin
    if(latches_23_write_sample) begin
      latches_23_storage = latches_23_write_data;
    end
  end

  assign latches_24_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h19)),(io_writes_0_valid && (io_writes_0_address == 6'h19))};
  assign latches_24_write_data = ((latches_24_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_24_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_24_write_sample = ((! clk) && latches_24_write_validReg);
  always @(*) begin
    if(latches_24_write_sample) begin
      latches_24_storage = latches_24_write_data;
    end
  end

  assign latches_25_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h1a)),(io_writes_0_valid && (io_writes_0_address == 6'h1a))};
  assign latches_25_write_data = ((latches_25_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_25_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_25_write_sample = ((! clk) && latches_25_write_validReg);
  always @(*) begin
    if(latches_25_write_sample) begin
      latches_25_storage = latches_25_write_data;
    end
  end

  assign latches_26_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h1b)),(io_writes_0_valid && (io_writes_0_address == 6'h1b))};
  assign latches_26_write_data = ((latches_26_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_26_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_26_write_sample = ((! clk) && latches_26_write_validReg);
  always @(*) begin
    if(latches_26_write_sample) begin
      latches_26_storage = latches_26_write_data;
    end
  end

  assign latches_27_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h1c)),(io_writes_0_valid && (io_writes_0_address == 6'h1c))};
  assign latches_27_write_data = ((latches_27_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_27_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_27_write_sample = ((! clk) && latches_27_write_validReg);
  always @(*) begin
    if(latches_27_write_sample) begin
      latches_27_storage = latches_27_write_data;
    end
  end

  assign latches_28_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h1d)),(io_writes_0_valid && (io_writes_0_address == 6'h1d))};
  assign latches_28_write_data = ((latches_28_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_28_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_28_write_sample = ((! clk) && latches_28_write_validReg);
  always @(*) begin
    if(latches_28_write_sample) begin
      latches_28_storage = latches_28_write_data;
    end
  end

  assign latches_29_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h1e)),(io_writes_0_valid && (io_writes_0_address == 6'h1e))};
  assign latches_29_write_data = ((latches_29_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_29_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_29_write_sample = ((! clk) && latches_29_write_validReg);
  always @(*) begin
    if(latches_29_write_sample) begin
      latches_29_storage = latches_29_write_data;
    end
  end

  assign latches_30_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h1f)),(io_writes_0_valid && (io_writes_0_address == 6'h1f))};
  assign latches_30_write_data = ((latches_30_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_30_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_30_write_sample = ((! clk) && latches_30_write_validReg);
  always @(*) begin
    if(latches_30_write_sample) begin
      latches_30_storage = latches_30_write_data;
    end
  end

  assign latches_31_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h20)),(io_writes_0_valid && (io_writes_0_address == 6'h20))};
  assign latches_31_write_data = ((latches_31_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_31_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_31_write_sample = ((! clk) && latches_31_write_validReg);
  always @(*) begin
    if(latches_31_write_sample) begin
      latches_31_storage = latches_31_write_data;
    end
  end

  assign latches_32_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h21)),(io_writes_0_valid && (io_writes_0_address == 6'h21))};
  assign latches_32_write_data = ((latches_32_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_32_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_32_write_sample = ((! clk) && latches_32_write_validReg);
  always @(*) begin
    if(latches_32_write_sample) begin
      latches_32_storage = latches_32_write_data;
    end
  end

  assign latches_33_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h22)),(io_writes_0_valid && (io_writes_0_address == 6'h22))};
  assign latches_33_write_data = ((latches_33_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_33_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_33_write_sample = ((! clk) && latches_33_write_validReg);
  always @(*) begin
    if(latches_33_write_sample) begin
      latches_33_storage = latches_33_write_data;
    end
  end

  assign latches_34_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h23)),(io_writes_0_valid && (io_writes_0_address == 6'h23))};
  assign latches_34_write_data = ((latches_34_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_34_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_34_write_sample = ((! clk) && latches_34_write_validReg);
  always @(*) begin
    if(latches_34_write_sample) begin
      latches_34_storage = latches_34_write_data;
    end
  end

  assign latches_35_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h24)),(io_writes_0_valid && (io_writes_0_address == 6'h24))};
  assign latches_35_write_data = ((latches_35_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_35_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_35_write_sample = ((! clk) && latches_35_write_validReg);
  always @(*) begin
    if(latches_35_write_sample) begin
      latches_35_storage = latches_35_write_data;
    end
  end

  assign latches_36_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h25)),(io_writes_0_valid && (io_writes_0_address == 6'h25))};
  assign latches_36_write_data = ((latches_36_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_36_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_36_write_sample = ((! clk) && latches_36_write_validReg);
  always @(*) begin
    if(latches_36_write_sample) begin
      latches_36_storage = latches_36_write_data;
    end
  end

  assign latches_37_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h26)),(io_writes_0_valid && (io_writes_0_address == 6'h26))};
  assign latches_37_write_data = ((latches_37_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_37_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_37_write_sample = ((! clk) && latches_37_write_validReg);
  always @(*) begin
    if(latches_37_write_sample) begin
      latches_37_storage = latches_37_write_data;
    end
  end

  assign latches_38_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h27)),(io_writes_0_valid && (io_writes_0_address == 6'h27))};
  assign latches_38_write_data = ((latches_38_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_38_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_38_write_sample = ((! clk) && latches_38_write_validReg);
  always @(*) begin
    if(latches_38_write_sample) begin
      latches_38_storage = latches_38_write_data;
    end
  end

  assign latches_39_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h28)),(io_writes_0_valid && (io_writes_0_address == 6'h28))};
  assign latches_39_write_data = ((latches_39_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_39_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_39_write_sample = ((! clk) && latches_39_write_validReg);
  always @(*) begin
    if(latches_39_write_sample) begin
      latches_39_storage = latches_39_write_data;
    end
  end

  assign latches_40_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h29)),(io_writes_0_valid && (io_writes_0_address == 6'h29))};
  assign latches_40_write_data = ((latches_40_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_40_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_40_write_sample = ((! clk) && latches_40_write_validReg);
  always @(*) begin
    if(latches_40_write_sample) begin
      latches_40_storage = latches_40_write_data;
    end
  end

  assign latches_41_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h2a)),(io_writes_0_valid && (io_writes_0_address == 6'h2a))};
  assign latches_41_write_data = ((latches_41_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_41_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_41_write_sample = ((! clk) && latches_41_write_validReg);
  always @(*) begin
    if(latches_41_write_sample) begin
      latches_41_storage = latches_41_write_data;
    end
  end

  assign latches_42_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h2b)),(io_writes_0_valid && (io_writes_0_address == 6'h2b))};
  assign latches_42_write_data = ((latches_42_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_42_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_42_write_sample = ((! clk) && latches_42_write_validReg);
  always @(*) begin
    if(latches_42_write_sample) begin
      latches_42_storage = latches_42_write_data;
    end
  end

  assign latches_43_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h2c)),(io_writes_0_valid && (io_writes_0_address == 6'h2c))};
  assign latches_43_write_data = ((latches_43_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_43_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_43_write_sample = ((! clk) && latches_43_write_validReg);
  always @(*) begin
    if(latches_43_write_sample) begin
      latches_43_storage = latches_43_write_data;
    end
  end

  assign latches_44_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h2d)),(io_writes_0_valid && (io_writes_0_address == 6'h2d))};
  assign latches_44_write_data = ((latches_44_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_44_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_44_write_sample = ((! clk) && latches_44_write_validReg);
  always @(*) begin
    if(latches_44_write_sample) begin
      latches_44_storage = latches_44_write_data;
    end
  end

  assign latches_45_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h2e)),(io_writes_0_valid && (io_writes_0_address == 6'h2e))};
  assign latches_45_write_data = ((latches_45_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_45_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_45_write_sample = ((! clk) && latches_45_write_validReg);
  always @(*) begin
    if(latches_45_write_sample) begin
      latches_45_storage = latches_45_write_data;
    end
  end

  assign latches_46_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h2f)),(io_writes_0_valid && (io_writes_0_address == 6'h2f))};
  assign latches_46_write_data = ((latches_46_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_46_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_46_write_sample = ((! clk) && latches_46_write_validReg);
  always @(*) begin
    if(latches_46_write_sample) begin
      latches_46_storage = latches_46_write_data;
    end
  end

  assign latches_47_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h30)),(io_writes_0_valid && (io_writes_0_address == 6'h30))};
  assign latches_47_write_data = ((latches_47_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_47_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_47_write_sample = ((! clk) && latches_47_write_validReg);
  always @(*) begin
    if(latches_47_write_sample) begin
      latches_47_storage = latches_47_write_data;
    end
  end

  assign latches_48_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h31)),(io_writes_0_valid && (io_writes_0_address == 6'h31))};
  assign latches_48_write_data = ((latches_48_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_48_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_48_write_sample = ((! clk) && latches_48_write_validReg);
  always @(*) begin
    if(latches_48_write_sample) begin
      latches_48_storage = latches_48_write_data;
    end
  end

  assign latches_49_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h32)),(io_writes_0_valid && (io_writes_0_address == 6'h32))};
  assign latches_49_write_data = ((latches_49_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_49_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_49_write_sample = ((! clk) && latches_49_write_validReg);
  always @(*) begin
    if(latches_49_write_sample) begin
      latches_49_storage = latches_49_write_data;
    end
  end

  assign latches_50_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h33)),(io_writes_0_valid && (io_writes_0_address == 6'h33))};
  assign latches_50_write_data = ((latches_50_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_50_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_50_write_sample = ((! clk) && latches_50_write_validReg);
  always @(*) begin
    if(latches_50_write_sample) begin
      latches_50_storage = latches_50_write_data;
    end
  end

  assign latches_51_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h34)),(io_writes_0_valid && (io_writes_0_address == 6'h34))};
  assign latches_51_write_data = ((latches_51_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_51_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_51_write_sample = ((! clk) && latches_51_write_validReg);
  always @(*) begin
    if(latches_51_write_sample) begin
      latches_51_storage = latches_51_write_data;
    end
  end

  assign latches_52_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h35)),(io_writes_0_valid && (io_writes_0_address == 6'h35))};
  assign latches_52_write_data = ((latches_52_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_52_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_52_write_sample = ((! clk) && latches_52_write_validReg);
  always @(*) begin
    if(latches_52_write_sample) begin
      latches_52_storage = latches_52_write_data;
    end
  end

  assign latches_53_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h36)),(io_writes_0_valid && (io_writes_0_address == 6'h36))};
  assign latches_53_write_data = ((latches_53_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_53_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_53_write_sample = ((! clk) && latches_53_write_validReg);
  always @(*) begin
    if(latches_53_write_sample) begin
      latches_53_storage = latches_53_write_data;
    end
  end

  assign latches_54_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h37)),(io_writes_0_valid && (io_writes_0_address == 6'h37))};
  assign latches_54_write_data = ((latches_54_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_54_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_54_write_sample = ((! clk) && latches_54_write_validReg);
  always @(*) begin
    if(latches_54_write_sample) begin
      latches_54_storage = latches_54_write_data;
    end
  end

  assign latches_55_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h38)),(io_writes_0_valid && (io_writes_0_address == 6'h38))};
  assign latches_55_write_data = ((latches_55_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_55_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_55_write_sample = ((! clk) && latches_55_write_validReg);
  always @(*) begin
    if(latches_55_write_sample) begin
      latches_55_storage = latches_55_write_data;
    end
  end

  assign latches_56_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h39)),(io_writes_0_valid && (io_writes_0_address == 6'h39))};
  assign latches_56_write_data = ((latches_56_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_56_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_56_write_sample = ((! clk) && latches_56_write_validReg);
  always @(*) begin
    if(latches_56_write_sample) begin
      latches_56_storage = latches_56_write_data;
    end
  end

  assign latches_57_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h3a)),(io_writes_0_valid && (io_writes_0_address == 6'h3a))};
  assign latches_57_write_data = ((latches_57_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_57_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_57_write_sample = ((! clk) && latches_57_write_validReg);
  always @(*) begin
    if(latches_57_write_sample) begin
      latches_57_storage = latches_57_write_data;
    end
  end

  assign latches_58_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h3b)),(io_writes_0_valid && (io_writes_0_address == 6'h3b))};
  assign latches_58_write_data = ((latches_58_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_58_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_58_write_sample = ((! clk) && latches_58_write_validReg);
  always @(*) begin
    if(latches_58_write_sample) begin
      latches_58_storage = latches_58_write_data;
    end
  end

  assign latches_59_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h3c)),(io_writes_0_valid && (io_writes_0_address == 6'h3c))};
  assign latches_59_write_data = ((latches_59_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_59_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_59_write_sample = ((! clk) && latches_59_write_validReg);
  always @(*) begin
    if(latches_59_write_sample) begin
      latches_59_storage = latches_59_write_data;
    end
  end

  assign latches_60_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h3d)),(io_writes_0_valid && (io_writes_0_address == 6'h3d))};
  assign latches_60_write_data = ((latches_60_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_60_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_60_write_sample = ((! clk) && latches_60_write_validReg);
  always @(*) begin
    if(latches_60_write_sample) begin
      latches_60_storage = latches_60_write_data;
    end
  end

  assign latches_61_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h3e)),(io_writes_0_valid && (io_writes_0_address == 6'h3e))};
  assign latches_61_write_data = ((latches_61_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_61_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_61_write_sample = ((! clk) && latches_61_write_validReg);
  always @(*) begin
    if(latches_61_write_sample) begin
      latches_61_storage = latches_61_write_data;
    end
  end

  assign latches_62_write_mask = {(io_writes_1_valid && (io_writes_1_address == 6'h3f)),(io_writes_0_valid && (io_writes_0_address == 6'h3f))};
  assign latches_62_write_data = ((latches_62_write_maskReg[0] ? writeFrontend_buffers_0 : 32'h00000000) | (latches_62_write_maskReg[1] ? writeFrontend_buffers_1 : 32'h00000000));
  assign latches_62_write_sample = ((! clk) && latches_62_write_validReg);
  always @(*) begin
    if(latches_62_write_sample) begin
      latches_62_storage = latches_62_write_data;
    end
  end

  assign readLogic_0_oh = (64'h0000000000000001 <<< io_reads_0_address);
  assign _zz_1 = readLogic_0_oh;
  assign io_reads_0_data = readLogic_0_tri;
  assign readLogic_1_oh = (64'h0000000000000001 <<< io_reads_1_address);
  assign _zz_2 = readLogic_1_oh;
  assign io_reads_1_data = readLogic_1_tri;
  assign readLogic_2_oh = (64'h0000000000000001 <<< io_reads_2_address);
  assign _zz_3 = readLogic_2_oh;
  assign io_reads_2_data = readLogic_2_tri;
  assign readLogic_3_oh = (64'h0000000000000001 <<< io_reads_3_address);
  assign _zz_4 = readLogic_3_oh;
  assign io_reads_3_data = readLogic_3_tri;
  always @(posedge clk) begin
    writeFrontend_buffers_0 <= io_writes_0_data;
    writeFrontend_buffers_1 <= io_writes_1_data;
    latches_0_write_maskReg <= latches_0_write_mask;
    latches_0_write_validReg <= (|latches_0_write_mask);
    latches_1_write_maskReg <= latches_1_write_mask;
    latches_1_write_validReg <= (|latches_1_write_mask);
    latches_2_write_maskReg <= latches_2_write_mask;
    latches_2_write_validReg <= (|latches_2_write_mask);
    latches_3_write_maskReg <= latches_3_write_mask;
    latches_3_write_validReg <= (|latches_3_write_mask);
    latches_4_write_maskReg <= latches_4_write_mask;
    latches_4_write_validReg <= (|latches_4_write_mask);
    latches_5_write_maskReg <= latches_5_write_mask;
    latches_5_write_validReg <= (|latches_5_write_mask);
    latches_6_write_maskReg <= latches_6_write_mask;
    latches_6_write_validReg <= (|latches_6_write_mask);
    latches_7_write_maskReg <= latches_7_write_mask;
    latches_7_write_validReg <= (|latches_7_write_mask);
    latches_8_write_maskReg <= latches_8_write_mask;
    latches_8_write_validReg <= (|latches_8_write_mask);
    latches_9_write_maskReg <= latches_9_write_mask;
    latches_9_write_validReg <= (|latches_9_write_mask);
    latches_10_write_maskReg <= latches_10_write_mask;
    latches_10_write_validReg <= (|latches_10_write_mask);
    latches_11_write_maskReg <= latches_11_write_mask;
    latches_11_write_validReg <= (|latches_11_write_mask);
    latches_12_write_maskReg <= latches_12_write_mask;
    latches_12_write_validReg <= (|latches_12_write_mask);
    latches_13_write_maskReg <= latches_13_write_mask;
    latches_13_write_validReg <= (|latches_13_write_mask);
    latches_14_write_maskReg <= latches_14_write_mask;
    latches_14_write_validReg <= (|latches_14_write_mask);
    latches_15_write_maskReg <= latches_15_write_mask;
    latches_15_write_validReg <= (|latches_15_write_mask);
    latches_16_write_maskReg <= latches_16_write_mask;
    latches_16_write_validReg <= (|latches_16_write_mask);
    latches_17_write_maskReg <= latches_17_write_mask;
    latches_17_write_validReg <= (|latches_17_write_mask);
    latches_18_write_maskReg <= latches_18_write_mask;
    latches_18_write_validReg <= (|latches_18_write_mask);
    latches_19_write_maskReg <= latches_19_write_mask;
    latches_19_write_validReg <= (|latches_19_write_mask);
    latches_20_write_maskReg <= latches_20_write_mask;
    latches_20_write_validReg <= (|latches_20_write_mask);
    latches_21_write_maskReg <= latches_21_write_mask;
    latches_21_write_validReg <= (|latches_21_write_mask);
    latches_22_write_maskReg <= latches_22_write_mask;
    latches_22_write_validReg <= (|latches_22_write_mask);
    latches_23_write_maskReg <= latches_23_write_mask;
    latches_23_write_validReg <= (|latches_23_write_mask);
    latches_24_write_maskReg <= latches_24_write_mask;
    latches_24_write_validReg <= (|latches_24_write_mask);
    latches_25_write_maskReg <= latches_25_write_mask;
    latches_25_write_validReg <= (|latches_25_write_mask);
    latches_26_write_maskReg <= latches_26_write_mask;
    latches_26_write_validReg <= (|latches_26_write_mask);
    latches_27_write_maskReg <= latches_27_write_mask;
    latches_27_write_validReg <= (|latches_27_write_mask);
    latches_28_write_maskReg <= latches_28_write_mask;
    latches_28_write_validReg <= (|latches_28_write_mask);
    latches_29_write_maskReg <= latches_29_write_mask;
    latches_29_write_validReg <= (|latches_29_write_mask);
    latches_30_write_maskReg <= latches_30_write_mask;
    latches_30_write_validReg <= (|latches_30_write_mask);
    latches_31_write_maskReg <= latches_31_write_mask;
    latches_31_write_validReg <= (|latches_31_write_mask);
    latches_32_write_maskReg <= latches_32_write_mask;
    latches_32_write_validReg <= (|latches_32_write_mask);
    latches_33_write_maskReg <= latches_33_write_mask;
    latches_33_write_validReg <= (|latches_33_write_mask);
    latches_34_write_maskReg <= latches_34_write_mask;
    latches_34_write_validReg <= (|latches_34_write_mask);
    latches_35_write_maskReg <= latches_35_write_mask;
    latches_35_write_validReg <= (|latches_35_write_mask);
    latches_36_write_maskReg <= latches_36_write_mask;
    latches_36_write_validReg <= (|latches_36_write_mask);
    latches_37_write_maskReg <= latches_37_write_mask;
    latches_37_write_validReg <= (|latches_37_write_mask);
    latches_38_write_maskReg <= latches_38_write_mask;
    latches_38_write_validReg <= (|latches_38_write_mask);
    latches_39_write_maskReg <= latches_39_write_mask;
    latches_39_write_validReg <= (|latches_39_write_mask);
    latches_40_write_maskReg <= latches_40_write_mask;
    latches_40_write_validReg <= (|latches_40_write_mask);
    latches_41_write_maskReg <= latches_41_write_mask;
    latches_41_write_validReg <= (|latches_41_write_mask);
    latches_42_write_maskReg <= latches_42_write_mask;
    latches_42_write_validReg <= (|latches_42_write_mask);
    latches_43_write_maskReg <= latches_43_write_mask;
    latches_43_write_validReg <= (|latches_43_write_mask);
    latches_44_write_maskReg <= latches_44_write_mask;
    latches_44_write_validReg <= (|latches_44_write_mask);
    latches_45_write_maskReg <= latches_45_write_mask;
    latches_45_write_validReg <= (|latches_45_write_mask);
    latches_46_write_maskReg <= latches_46_write_mask;
    latches_46_write_validReg <= (|latches_46_write_mask);
    latches_47_write_maskReg <= latches_47_write_mask;
    latches_47_write_validReg <= (|latches_47_write_mask);
    latches_48_write_maskReg <= latches_48_write_mask;
    latches_48_write_validReg <= (|latches_48_write_mask);
    latches_49_write_maskReg <= latches_49_write_mask;
    latches_49_write_validReg <= (|latches_49_write_mask);
    latches_50_write_maskReg <= latches_50_write_mask;
    latches_50_write_validReg <= (|latches_50_write_mask);
    latches_51_write_maskReg <= latches_51_write_mask;
    latches_51_write_validReg <= (|latches_51_write_mask);
    latches_52_write_maskReg <= latches_52_write_mask;
    latches_52_write_validReg <= (|latches_52_write_mask);
    latches_53_write_maskReg <= latches_53_write_mask;
    latches_53_write_validReg <= (|latches_53_write_mask);
    latches_54_write_maskReg <= latches_54_write_mask;
    latches_54_write_validReg <= (|latches_54_write_mask);
    latches_55_write_maskReg <= latches_55_write_mask;
    latches_55_write_validReg <= (|latches_55_write_mask);
    latches_56_write_maskReg <= latches_56_write_mask;
    latches_56_write_validReg <= (|latches_56_write_mask);
    latches_57_write_maskReg <= latches_57_write_mask;
    latches_57_write_validReg <= (|latches_57_write_mask);
    latches_58_write_maskReg <= latches_58_write_mask;
    latches_58_write_validReg <= (|latches_58_write_mask);
    latches_59_write_maskReg <= latches_59_write_mask;
    latches_59_write_validReg <= (|latches_59_write_mask);
    latches_60_write_maskReg <= latches_60_write_mask;
    latches_60_write_validReg <= (|latches_60_write_mask);
    latches_61_write_maskReg <= latches_61_write_mask;
    latches_61_write_validReg <= (|latches_61_write_mask);
    latches_62_write_maskReg <= latches_62_write_mask;
    latches_62_write_validReg <= (|latches_62_write_mask);
  end


endmodule

module IssueQueue (
  input  wire          io_clear,
  (* keep , syn_keep *) input  wire [7:0]    io_events /* synthesis syn_keep = 1 */ ,
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [7:0]    io_push_payload_slots_0_event,
  input  wire [1:0]    io_push_payload_slots_0_sel,
  input  wire [0:0]    io_push_payload_slots_0_context_staticWake,
  input  wire [5:0]    io_push_payload_slots_0_context_physRd,
  input  wire [3:0]    io_push_payload_slots_0_context_robId,
  input  wire [5:0]    io_push_payload_slots_0_context_euCtx_0,
  input  wire [5:0]    io_push_payload_slots_0_context_euCtx_1,
  output wire          io_schedules_0_valid,
  input  wire          io_schedules_0_ready,
  output wire [7:0]    io_schedules_0_payload_event,
  output wire          io_schedules_1_valid,
  input  wire          io_schedules_1_ready,
  output wire [7:0]    io_schedules_1_payload_event,
  output wire [0:0]    io_contexts_0_staticWake,
  output wire [5:0]    io_contexts_0_physRd,
  output wire [3:0]    io_contexts_0_robId,
  output wire [5:0]    io_contexts_0_euCtx_0,
  output wire [5:0]    io_contexts_0_euCtx_1,
  output wire [0:0]    io_contexts_1_staticWake,
  output wire [5:0]    io_contexts_1_physRd,
  output wire [3:0]    io_contexts_1_robId,
  output wire [5:0]    io_contexts_1_euCtx_0,
  output wire [5:0]    io_contexts_1_euCtx_1,
  output wire [0:0]    io_contexts_2_staticWake,
  output wire [5:0]    io_contexts_2_physRd,
  output wire [3:0]    io_contexts_2_robId,
  output wire [5:0]    io_contexts_2_euCtx_0,
  output wire [5:0]    io_contexts_2_euCtx_1,
  output wire [0:0]    io_contexts_3_staticWake,
  output wire [5:0]    io_contexts_3_physRd,
  output wire [3:0]    io_contexts_3_robId,
  output wire [5:0]    io_contexts_3_euCtx_0,
  output wire [5:0]    io_contexts_3_euCtx_1,
  output wire [0:0]    io_contexts_4_staticWake,
  output wire [5:0]    io_contexts_4_physRd,
  output wire [3:0]    io_contexts_4_robId,
  output wire [5:0]    io_contexts_4_euCtx_0,
  output wire [5:0]    io_contexts_4_euCtx_1,
  output wire [0:0]    io_contexts_5_staticWake,
  output wire [5:0]    io_contexts_5_physRd,
  output wire [3:0]    io_contexts_5_robId,
  output wire [5:0]    io_contexts_5_euCtx_0,
  output wire [5:0]    io_contexts_5_euCtx_1,
  output wire [0:0]    io_contexts_6_staticWake,
  output wire [5:0]    io_contexts_6_physRd,
  output wire [3:0]    io_contexts_6_robId,
  output wire [5:0]    io_contexts_6_euCtx_0,
  output wire [5:0]    io_contexts_6_euCtx_1,
  output wire [0:0]    io_contexts_7_staticWake,
  output wire [5:0]    io_contexts_7_physRd,
  output wire [3:0]    io_contexts_7_robId,
  output wire [5:0]    io_contexts_7_euCtx_0,
  output wire [5:0]    io_contexts_7_euCtx_1,
  output reg  [7:0]    io_usage,
  input  wire          clk,
  input  wire          reset
);

  wire       [7:0]    _zz_event_moved;
  wire                _zz_selector_0_slotsValid;
  wire                _zz_selector_0_slotsValid_1;
  wire       [0:0]    _zz_selector_0_slotsValid_2;
  wire       [0:0]    _zz_selector_0_slotsValid_3;
  wire                _zz_selector_1_slotsValid;
  wire                _zz_selector_1_slotsValid_1;
  wire       [0:0]    _zz_selector_1_slotsValid_2;
  wire       [0:0]    _zz_selector_1_slotsValid_3;
  reg                 running;
  wire                clear;
  wire                lines_0_ways_0_fire;
  reg        [1:0]    lines_0_ways_0_sel;
  reg        [1:0]    lines_0_ways_0_selComb;
  reg        [0:0]    lines_0_ways_0_triggers;
  wire                lines_0_ways_0_ready;
  reg        [0:0]    lines_0_ways_0_context_staticWake;
  reg        [5:0]    lines_0_ways_0_context_physRd;
  reg        [3:0]    lines_0_ways_0_context_robId;
  reg        [5:0]    lines_0_ways_0_context_euCtx_0;
  reg        [5:0]    lines_0_ways_0_context_euCtx_1;
  wire                lines_1_ways_0_fire;
  reg        [1:0]    lines_1_ways_0_sel;
  reg        [1:0]    lines_1_ways_0_selComb;
  reg        [1:0]    lines_1_ways_0_triggers;
  wire                lines_1_ways_0_ready;
  reg        [0:0]    lines_1_ways_0_context_staticWake;
  reg        [5:0]    lines_1_ways_0_context_physRd;
  reg        [3:0]    lines_1_ways_0_context_robId;
  reg        [5:0]    lines_1_ways_0_context_euCtx_0;
  reg        [5:0]    lines_1_ways_0_context_euCtx_1;
  wire                lines_2_ways_0_fire;
  reg        [1:0]    lines_2_ways_0_sel;
  reg        [1:0]    lines_2_ways_0_selComb;
  reg        [2:0]    lines_2_ways_0_triggers;
  wire                lines_2_ways_0_ready;
  reg        [0:0]    lines_2_ways_0_context_staticWake;
  reg        [5:0]    lines_2_ways_0_context_physRd;
  reg        [3:0]    lines_2_ways_0_context_robId;
  reg        [5:0]    lines_2_ways_0_context_euCtx_0;
  reg        [5:0]    lines_2_ways_0_context_euCtx_1;
  wire                lines_3_ways_0_fire;
  reg        [1:0]    lines_3_ways_0_sel;
  reg        [1:0]    lines_3_ways_0_selComb;
  reg        [3:0]    lines_3_ways_0_triggers;
  wire                lines_3_ways_0_ready;
  reg        [0:0]    lines_3_ways_0_context_staticWake;
  reg        [5:0]    lines_3_ways_0_context_physRd;
  reg        [3:0]    lines_3_ways_0_context_robId;
  reg        [5:0]    lines_3_ways_0_context_euCtx_0;
  reg        [5:0]    lines_3_ways_0_context_euCtx_1;
  wire                lines_4_ways_0_fire;
  reg        [1:0]    lines_4_ways_0_sel;
  reg        [1:0]    lines_4_ways_0_selComb;
  reg        [4:0]    lines_4_ways_0_triggers;
  wire                lines_4_ways_0_ready;
  reg        [0:0]    lines_4_ways_0_context_staticWake;
  reg        [5:0]    lines_4_ways_0_context_physRd;
  reg        [3:0]    lines_4_ways_0_context_robId;
  reg        [5:0]    lines_4_ways_0_context_euCtx_0;
  reg        [5:0]    lines_4_ways_0_context_euCtx_1;
  wire                lines_5_ways_0_fire;
  reg        [1:0]    lines_5_ways_0_sel;
  reg        [1:0]    lines_5_ways_0_selComb;
  reg        [5:0]    lines_5_ways_0_triggers;
  wire                lines_5_ways_0_ready;
  reg        [0:0]    lines_5_ways_0_context_staticWake;
  reg        [5:0]    lines_5_ways_0_context_physRd;
  reg        [3:0]    lines_5_ways_0_context_robId;
  reg        [5:0]    lines_5_ways_0_context_euCtx_0;
  reg        [5:0]    lines_5_ways_0_context_euCtx_1;
  wire                lines_6_ways_0_fire;
  reg        [1:0]    lines_6_ways_0_sel;
  reg        [1:0]    lines_6_ways_0_selComb;
  reg        [6:0]    lines_6_ways_0_triggers;
  wire                lines_6_ways_0_ready;
  reg        [0:0]    lines_6_ways_0_context_staticWake;
  reg        [5:0]    lines_6_ways_0_context_physRd;
  reg        [3:0]    lines_6_ways_0_context_robId;
  reg        [5:0]    lines_6_ways_0_context_euCtx_0;
  reg        [5:0]    lines_6_ways_0_context_euCtx_1;
  wire                lines_7_ways_0_fire;
  reg        [1:0]    lines_7_ways_0_sel;
  reg        [1:0]    lines_7_ways_0_selComb;
  reg        [7:0]    lines_7_ways_0_triggers;
  wire                lines_7_ways_0_ready;
  reg        [0:0]    lines_7_ways_0_context_staticWake;
  reg        [5:0]    lines_7_ways_0_context_physRd;
  reg        [3:0]    lines_7_ways_0_context_robId;
  reg        [5:0]    lines_7_ways_0_context_euCtx_0;
  reg        [5:0]    lines_7_ways_0_context_euCtx_1;
  wire                compaction_moveIt;
  wire       [7:0]    event_moved;
  wire       [7:0]    event_value;
  wire                when_IssueQueue_l109;
  wire                when_IssueQueue_l109_1;
  wire                when_IssueQueue_l109_2;
  wire                when_IssueQueue_l109_3;
  wire                when_IssueQueue_l109_4;
  wire                when_IssueQueue_l109_5;
  wire                when_IssueQueue_l109_6;
  wire                when_IssueQueue_l109_7;
  wire       [7:0]    selector_0_slotsValid;
  wire       [7:0]    _zz_selector_0_slotsValid_bools_0;
  wire                selector_0_slotsValid_bools_0;
  wire                selector_0_slotsValid_bools_1;
  wire                selector_0_slotsValid_bools_2;
  wire                selector_0_slotsValid_bools_3;
  wire                selector_0_slotsValid_bools_4;
  wire                selector_0_slotsValid_bools_5;
  wire                selector_0_slotsValid_bools_6;
  wire                selector_0_slotsValid_bools_7;
  reg        [7:0]    _zz_selector_0_selOh;
  wire                selector_0_slotsValid_range_0_to_1;
  wire                selector_0_slotsValid_range_0_to_2;
  wire                selector_0_slotsValid_range_0_to_3;
  wire                selector_0_slotsValid_range_4_to_5;
  wire                selector_0_slotsValid_range_4_to_6;
  wire       [7:0]    selector_0_selOh;
  wire       [7:0]    selector_1_slotsValid;
  wire       [7:0]    _zz_selector_1_slotsValid_bools_0;
  wire                selector_1_slotsValid_bools_0;
  wire                selector_1_slotsValid_bools_1;
  wire                selector_1_slotsValid_bools_2;
  wire                selector_1_slotsValid_bools_3;
  wire                selector_1_slotsValid_bools_4;
  wire                selector_1_slotsValid_bools_5;
  wire                selector_1_slotsValid_bools_6;
  wire                selector_1_slotsValid_bools_7;
  reg        [7:0]    _zz_selector_1_selOh;
  wire                selector_1_slotsValid_range_0_to_1;
  wire                selector_1_slotsValid_range_0_to_2;
  wire                selector_1_slotsValid_range_0_to_3;
  wire                selector_1_slotsValid_range_4_to_5;
  wire                selector_1_slotsValid_range_4_to_6;
  wire       [7:0]    selector_1_selOh;
  wire                line0Ready;
  wire                line1Ready;
  reg                 readyReg;

  assign _zz_event_moved = (io_events >>> 1);
  assign _zz_selector_0_slotsValid = lines_3_ways_0_sel[0];
  assign _zz_selector_0_slotsValid_1 = (lines_2_ways_0_ready && lines_2_ways_0_sel[0]);
  assign _zz_selector_0_slotsValid_2 = (lines_1_ways_0_ready && lines_1_ways_0_sel[0]);
  assign _zz_selector_0_slotsValid_3 = (lines_0_ways_0_ready && lines_0_ways_0_sel[0]);
  assign _zz_selector_1_slotsValid = lines_3_ways_0_sel[1];
  assign _zz_selector_1_slotsValid_1 = (lines_2_ways_0_ready && lines_2_ways_0_sel[1]);
  assign _zz_selector_1_slotsValid_2 = (lines_1_ways_0_ready && lines_1_ways_0_sel[1]);
  assign _zz_selector_1_slotsValid_3 = (lines_0_ways_0_ready && lines_0_ways_0_sel[1]);
  assign clear = (io_clear || (! running));
  always @(*) begin
    lines_0_ways_0_selComb = lines_0_ways_0_sel;
    if(lines_0_ways_0_fire) begin
      lines_0_ways_0_selComb = 2'b00;
    end
  end

  assign lines_0_ways_0_ready = 1'b1;
  assign io_contexts_0_staticWake = lines_0_ways_0_context_staticWake;
  assign io_contexts_0_physRd = lines_0_ways_0_context_physRd;
  assign io_contexts_0_robId = lines_0_ways_0_context_robId;
  assign io_contexts_0_euCtx_0 = lines_0_ways_0_context_euCtx_0;
  assign io_contexts_0_euCtx_1 = lines_0_ways_0_context_euCtx_1;
  always @(*) begin
    io_usage[0] = ((lines_0_ways_0_sel != 2'b00) || lines_0_ways_0_triggers[0]);
    io_usage[1] = ((lines_1_ways_0_sel != 2'b00) || lines_1_ways_0_triggers[1]);
    io_usage[2] = ((lines_2_ways_0_sel != 2'b00) || lines_2_ways_0_triggers[2]);
    io_usage[3] = ((lines_3_ways_0_sel != 2'b00) || lines_3_ways_0_triggers[3]);
    io_usage[4] = ((lines_4_ways_0_sel != 2'b00) || lines_4_ways_0_triggers[4]);
    io_usage[5] = ((lines_5_ways_0_sel != 2'b00) || lines_5_ways_0_triggers[5]);
    io_usage[6] = ((lines_6_ways_0_sel != 2'b00) || lines_6_ways_0_triggers[6]);
    io_usage[7] = ((lines_7_ways_0_sel != 2'b00) || lines_7_ways_0_triggers[7]);
  end

  always @(*) begin
    lines_1_ways_0_selComb = lines_1_ways_0_sel;
    if(lines_1_ways_0_fire) begin
      lines_1_ways_0_selComb = 2'b00;
    end
  end

  assign lines_1_ways_0_ready = (lines_1_ways_0_triggers[0 : 0] == 1'b0);
  assign io_contexts_1_staticWake = lines_1_ways_0_context_staticWake;
  assign io_contexts_1_physRd = lines_1_ways_0_context_physRd;
  assign io_contexts_1_robId = lines_1_ways_0_context_robId;
  assign io_contexts_1_euCtx_0 = lines_1_ways_0_context_euCtx_0;
  assign io_contexts_1_euCtx_1 = lines_1_ways_0_context_euCtx_1;
  always @(*) begin
    lines_2_ways_0_selComb = lines_2_ways_0_sel;
    if(lines_2_ways_0_fire) begin
      lines_2_ways_0_selComb = 2'b00;
    end
  end

  assign lines_2_ways_0_ready = (lines_2_ways_0_triggers[1 : 0] == 2'b00);
  assign io_contexts_2_staticWake = lines_2_ways_0_context_staticWake;
  assign io_contexts_2_physRd = lines_2_ways_0_context_physRd;
  assign io_contexts_2_robId = lines_2_ways_0_context_robId;
  assign io_contexts_2_euCtx_0 = lines_2_ways_0_context_euCtx_0;
  assign io_contexts_2_euCtx_1 = lines_2_ways_0_context_euCtx_1;
  always @(*) begin
    lines_3_ways_0_selComb = lines_3_ways_0_sel;
    if(lines_3_ways_0_fire) begin
      lines_3_ways_0_selComb = 2'b00;
    end
  end

  assign lines_3_ways_0_ready = (lines_3_ways_0_triggers[2 : 0] == 3'b000);
  assign io_contexts_3_staticWake = lines_3_ways_0_context_staticWake;
  assign io_contexts_3_physRd = lines_3_ways_0_context_physRd;
  assign io_contexts_3_robId = lines_3_ways_0_context_robId;
  assign io_contexts_3_euCtx_0 = lines_3_ways_0_context_euCtx_0;
  assign io_contexts_3_euCtx_1 = lines_3_ways_0_context_euCtx_1;
  always @(*) begin
    lines_4_ways_0_selComb = lines_4_ways_0_sel;
    if(lines_4_ways_0_fire) begin
      lines_4_ways_0_selComb = 2'b00;
    end
  end

  assign lines_4_ways_0_ready = (lines_4_ways_0_triggers[3 : 0] == 4'b0000);
  assign io_contexts_4_staticWake = lines_4_ways_0_context_staticWake;
  assign io_contexts_4_physRd = lines_4_ways_0_context_physRd;
  assign io_contexts_4_robId = lines_4_ways_0_context_robId;
  assign io_contexts_4_euCtx_0 = lines_4_ways_0_context_euCtx_0;
  assign io_contexts_4_euCtx_1 = lines_4_ways_0_context_euCtx_1;
  always @(*) begin
    lines_5_ways_0_selComb = lines_5_ways_0_sel;
    if(lines_5_ways_0_fire) begin
      lines_5_ways_0_selComb = 2'b00;
    end
  end

  assign lines_5_ways_0_ready = (lines_5_ways_0_triggers[4 : 0] == 5'h00);
  assign io_contexts_5_staticWake = lines_5_ways_0_context_staticWake;
  assign io_contexts_5_physRd = lines_5_ways_0_context_physRd;
  assign io_contexts_5_robId = lines_5_ways_0_context_robId;
  assign io_contexts_5_euCtx_0 = lines_5_ways_0_context_euCtx_0;
  assign io_contexts_5_euCtx_1 = lines_5_ways_0_context_euCtx_1;
  always @(*) begin
    lines_6_ways_0_selComb = lines_6_ways_0_sel;
    if(lines_6_ways_0_fire) begin
      lines_6_ways_0_selComb = 2'b00;
    end
  end

  assign lines_6_ways_0_ready = (lines_6_ways_0_triggers[5 : 0] == 6'h00);
  assign io_contexts_6_staticWake = lines_6_ways_0_context_staticWake;
  assign io_contexts_6_physRd = lines_6_ways_0_context_physRd;
  assign io_contexts_6_robId = lines_6_ways_0_context_robId;
  assign io_contexts_6_euCtx_0 = lines_6_ways_0_context_euCtx_0;
  assign io_contexts_6_euCtx_1 = lines_6_ways_0_context_euCtx_1;
  always @(*) begin
    lines_7_ways_0_selComb = lines_7_ways_0_sel;
    if(lines_7_ways_0_fire) begin
      lines_7_ways_0_selComb = 2'b00;
    end
  end

  assign lines_7_ways_0_ready = (lines_7_ways_0_triggers[6 : 0] == 7'h00);
  assign io_contexts_7_staticWake = lines_7_ways_0_context_staticWake;
  assign io_contexts_7_physRd = lines_7_ways_0_context_physRd;
  assign io_contexts_7_robId = lines_7_ways_0_context_robId;
  assign io_contexts_7_euCtx_0 = lines_7_ways_0_context_euCtx_0;
  assign io_contexts_7_euCtx_1 = lines_7_ways_0_context_euCtx_1;
  assign compaction_moveIt = (io_push_valid && io_push_ready);
  assign event_moved = ((! compaction_moveIt) ? io_events : _zz_event_moved);
  assign event_value = (clear ? 8'hff : event_moved);
  assign when_IssueQueue_l109 = event_value[0];
  assign when_IssueQueue_l109_1 = event_value[1];
  assign when_IssueQueue_l109_2 = event_value[2];
  assign when_IssueQueue_l109_3 = event_value[3];
  assign when_IssueQueue_l109_4 = event_value[4];
  assign when_IssueQueue_l109_5 = event_value[5];
  assign when_IssueQueue_l109_6 = event_value[6];
  assign when_IssueQueue_l109_7 = event_value[7];
  assign selector_0_slotsValid = {(lines_7_ways_0_ready && lines_7_ways_0_sel[0]),{(lines_6_ways_0_ready && lines_6_ways_0_sel[0]),{(lines_5_ways_0_ready && lines_5_ways_0_sel[0]),{(lines_4_ways_0_ready && lines_4_ways_0_sel[0]),{(lines_3_ways_0_ready && _zz_selector_0_slotsValid),{_zz_selector_0_slotsValid_1,{_zz_selector_0_slotsValid_2,_zz_selector_0_slotsValid_3}}}}}}};
  assign _zz_selector_0_slotsValid_bools_0 = selector_0_slotsValid;
  assign selector_0_slotsValid_bools_0 = _zz_selector_0_slotsValid_bools_0[0];
  assign selector_0_slotsValid_bools_1 = _zz_selector_0_slotsValid_bools_0[1];
  assign selector_0_slotsValid_bools_2 = _zz_selector_0_slotsValid_bools_0[2];
  assign selector_0_slotsValid_bools_3 = _zz_selector_0_slotsValid_bools_0[3];
  assign selector_0_slotsValid_bools_4 = _zz_selector_0_slotsValid_bools_0[4];
  assign selector_0_slotsValid_bools_5 = _zz_selector_0_slotsValid_bools_0[5];
  assign selector_0_slotsValid_bools_6 = _zz_selector_0_slotsValid_bools_0[6];
  assign selector_0_slotsValid_bools_7 = _zz_selector_0_slotsValid_bools_0[7];
  always @(*) begin
    _zz_selector_0_selOh[0] = (selector_0_slotsValid_bools_0 && (! 1'b0));
    _zz_selector_0_selOh[1] = (selector_0_slotsValid_bools_1 && (! selector_0_slotsValid_bools_0));
    _zz_selector_0_selOh[2] = (selector_0_slotsValid_bools_2 && (! selector_0_slotsValid_range_0_to_1));
    _zz_selector_0_selOh[3] = (selector_0_slotsValid_bools_3 && (! selector_0_slotsValid_range_0_to_2));
    _zz_selector_0_selOh[4] = (selector_0_slotsValid_bools_4 && (! selector_0_slotsValid_range_0_to_3));
    _zz_selector_0_selOh[5] = (selector_0_slotsValid_bools_5 && (! (selector_0_slotsValid_bools_4 || selector_0_slotsValid_range_0_to_3)));
    _zz_selector_0_selOh[6] = (selector_0_slotsValid_bools_6 && (! (selector_0_slotsValid_range_4_to_5 || selector_0_slotsValid_range_0_to_3)));
    _zz_selector_0_selOh[7] = (selector_0_slotsValid_bools_7 && (! (selector_0_slotsValid_range_4_to_6 || selector_0_slotsValid_range_0_to_3)));
  end

  assign selector_0_slotsValid_range_0_to_1 = (|{selector_0_slotsValid_bools_1,selector_0_slotsValid_bools_0});
  assign selector_0_slotsValid_range_0_to_2 = (|{selector_0_slotsValid_bools_2,{selector_0_slotsValid_bools_1,selector_0_slotsValid_bools_0}});
  assign selector_0_slotsValid_range_0_to_3 = (|{selector_0_slotsValid_bools_3,{selector_0_slotsValid_bools_2,{selector_0_slotsValid_bools_1,selector_0_slotsValid_bools_0}}});
  assign selector_0_slotsValid_range_4_to_5 = (|{selector_0_slotsValid_bools_5,selector_0_slotsValid_bools_4});
  assign selector_0_slotsValid_range_4_to_6 = (|{selector_0_slotsValid_bools_6,{selector_0_slotsValid_bools_5,selector_0_slotsValid_bools_4}});
  assign selector_0_selOh = _zz_selector_0_selOh;
  assign io_schedules_0_valid = ((|selector_0_slotsValid) && running);
  assign io_schedules_0_payload_event = selector_0_selOh;
  assign selector_1_slotsValid = {(lines_7_ways_0_ready && lines_7_ways_0_sel[1]),{(lines_6_ways_0_ready && lines_6_ways_0_sel[1]),{(lines_5_ways_0_ready && lines_5_ways_0_sel[1]),{(lines_4_ways_0_ready && lines_4_ways_0_sel[1]),{(lines_3_ways_0_ready && _zz_selector_1_slotsValid),{_zz_selector_1_slotsValid_1,{_zz_selector_1_slotsValid_2,_zz_selector_1_slotsValid_3}}}}}}};
  assign _zz_selector_1_slotsValid_bools_0 = selector_1_slotsValid;
  assign selector_1_slotsValid_bools_0 = _zz_selector_1_slotsValid_bools_0[0];
  assign selector_1_slotsValid_bools_1 = _zz_selector_1_slotsValid_bools_0[1];
  assign selector_1_slotsValid_bools_2 = _zz_selector_1_slotsValid_bools_0[2];
  assign selector_1_slotsValid_bools_3 = _zz_selector_1_slotsValid_bools_0[3];
  assign selector_1_slotsValid_bools_4 = _zz_selector_1_slotsValid_bools_0[4];
  assign selector_1_slotsValid_bools_5 = _zz_selector_1_slotsValid_bools_0[5];
  assign selector_1_slotsValid_bools_6 = _zz_selector_1_slotsValid_bools_0[6];
  assign selector_1_slotsValid_bools_7 = _zz_selector_1_slotsValid_bools_0[7];
  always @(*) begin
    _zz_selector_1_selOh[0] = (selector_1_slotsValid_bools_0 && (! 1'b0));
    _zz_selector_1_selOh[1] = (selector_1_slotsValid_bools_1 && (! selector_1_slotsValid_bools_0));
    _zz_selector_1_selOh[2] = (selector_1_slotsValid_bools_2 && (! selector_1_slotsValid_range_0_to_1));
    _zz_selector_1_selOh[3] = (selector_1_slotsValid_bools_3 && (! selector_1_slotsValid_range_0_to_2));
    _zz_selector_1_selOh[4] = (selector_1_slotsValid_bools_4 && (! selector_1_slotsValid_range_0_to_3));
    _zz_selector_1_selOh[5] = (selector_1_slotsValid_bools_5 && (! (selector_1_slotsValid_bools_4 || selector_1_slotsValid_range_0_to_3)));
    _zz_selector_1_selOh[6] = (selector_1_slotsValid_bools_6 && (! (selector_1_slotsValid_range_4_to_5 || selector_1_slotsValid_range_0_to_3)));
    _zz_selector_1_selOh[7] = (selector_1_slotsValid_bools_7 && (! (selector_1_slotsValid_range_4_to_6 || selector_1_slotsValid_range_0_to_3)));
  end

  assign selector_1_slotsValid_range_0_to_1 = (|{selector_1_slotsValid_bools_1,selector_1_slotsValid_bools_0});
  assign selector_1_slotsValid_range_0_to_2 = (|{selector_1_slotsValid_bools_2,{selector_1_slotsValid_bools_1,selector_1_slotsValid_bools_0}});
  assign selector_1_slotsValid_range_0_to_3 = (|{selector_1_slotsValid_bools_3,{selector_1_slotsValid_bools_2,{selector_1_slotsValid_bools_1,selector_1_slotsValid_bools_0}}});
  assign selector_1_slotsValid_range_4_to_5 = (|{selector_1_slotsValid_bools_5,selector_1_slotsValid_bools_4});
  assign selector_1_slotsValid_range_4_to_6 = (|{selector_1_slotsValid_bools_6,{selector_1_slotsValid_bools_5,selector_1_slotsValid_bools_4}});
  assign selector_1_selOh = _zz_selector_1_selOh;
  assign io_schedules_1_valid = ((|selector_1_slotsValid) && running);
  assign io_schedules_1_payload_event = selector_1_selOh;
  assign lines_0_ways_0_fire = (|{(io_schedules_1_ready && selector_1_selOh[0]),(io_schedules_0_ready && selector_0_selOh[0])});
  assign lines_1_ways_0_fire = (|{(io_schedules_1_ready && selector_1_selOh[1]),(io_schedules_0_ready && selector_0_selOh[1])});
  assign lines_2_ways_0_fire = (|{(io_schedules_1_ready && selector_1_selOh[2]),(io_schedules_0_ready && selector_0_selOh[2])});
  assign lines_3_ways_0_fire = (|{(io_schedules_1_ready && selector_1_selOh[3]),(io_schedules_0_ready && selector_0_selOh[3])});
  assign lines_4_ways_0_fire = (|{(io_schedules_1_ready && selector_1_selOh[4]),(io_schedules_0_ready && selector_0_selOh[4])});
  assign lines_5_ways_0_fire = (|{(io_schedules_1_ready && selector_1_selOh[5]),(io_schedules_0_ready && selector_0_selOh[5])});
  assign lines_6_ways_0_fire = (|{(io_schedules_1_ready && selector_1_selOh[6]),(io_schedules_0_ready && selector_0_selOh[6])});
  assign lines_7_ways_0_fire = (|{(io_schedules_1_ready && selector_1_selOh[7]),(io_schedules_0_ready && selector_0_selOh[7])});
  assign line0Ready = (&((! lines_0_ways_0_triggers[0]) && (lines_0_ways_0_sel == 2'b00)));
  assign line1Ready = (&((! lines_1_ways_0_triggers[1]) && (lines_1_ways_0_sel == 2'b00)));
  assign io_push_ready = readyReg;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      running <= 1'b0;
      readyReg <= 1'b0;
    end else begin
      running <= 1'b1;
      readyReg <= (compaction_moveIt ? line1Ready : line0Ready);
    end
  end

  always @(posedge clk) begin
    lines_0_ways_0_sel <= lines_0_ways_0_selComb;
    lines_1_ways_0_sel <= lines_1_ways_0_selComb;
    lines_2_ways_0_sel <= lines_2_ways_0_selComb;
    lines_3_ways_0_sel <= lines_3_ways_0_selComb;
    lines_4_ways_0_sel <= lines_4_ways_0_selComb;
    lines_5_ways_0_sel <= lines_5_ways_0_selComb;
    lines_6_ways_0_sel <= lines_6_ways_0_selComb;
    lines_7_ways_0_sel <= lines_7_ways_0_selComb;
    if(compaction_moveIt) begin
      lines_0_ways_0_context_staticWake <= lines_1_ways_0_context_staticWake;
      lines_0_ways_0_context_physRd <= lines_1_ways_0_context_physRd;
      lines_0_ways_0_context_robId <= lines_1_ways_0_context_robId;
      lines_0_ways_0_context_euCtx_0 <= lines_1_ways_0_context_euCtx_0;
      lines_0_ways_0_context_euCtx_1 <= lines_1_ways_0_context_euCtx_1;
      lines_0_ways_0_triggers <= (lines_1_ways_0_triggers >>> 1'd1);
      lines_0_ways_0_sel <= lines_1_ways_0_selComb;
      lines_1_ways_0_context_staticWake <= lines_2_ways_0_context_staticWake;
      lines_1_ways_0_context_physRd <= lines_2_ways_0_context_physRd;
      lines_1_ways_0_context_robId <= lines_2_ways_0_context_robId;
      lines_1_ways_0_context_euCtx_0 <= lines_2_ways_0_context_euCtx_0;
      lines_1_ways_0_context_euCtx_1 <= lines_2_ways_0_context_euCtx_1;
      lines_1_ways_0_triggers <= (lines_2_ways_0_triggers >>> 1'd1);
      lines_1_ways_0_sel <= lines_2_ways_0_selComb;
      lines_2_ways_0_context_staticWake <= lines_3_ways_0_context_staticWake;
      lines_2_ways_0_context_physRd <= lines_3_ways_0_context_physRd;
      lines_2_ways_0_context_robId <= lines_3_ways_0_context_robId;
      lines_2_ways_0_context_euCtx_0 <= lines_3_ways_0_context_euCtx_0;
      lines_2_ways_0_context_euCtx_1 <= lines_3_ways_0_context_euCtx_1;
      lines_2_ways_0_triggers <= (lines_3_ways_0_triggers >>> 1'd1);
      lines_2_ways_0_sel <= lines_3_ways_0_selComb;
      lines_3_ways_0_context_staticWake <= lines_4_ways_0_context_staticWake;
      lines_3_ways_0_context_physRd <= lines_4_ways_0_context_physRd;
      lines_3_ways_0_context_robId <= lines_4_ways_0_context_robId;
      lines_3_ways_0_context_euCtx_0 <= lines_4_ways_0_context_euCtx_0;
      lines_3_ways_0_context_euCtx_1 <= lines_4_ways_0_context_euCtx_1;
      lines_3_ways_0_triggers <= (lines_4_ways_0_triggers >>> 1'd1);
      lines_3_ways_0_sel <= lines_4_ways_0_selComb;
      lines_4_ways_0_context_staticWake <= lines_5_ways_0_context_staticWake;
      lines_4_ways_0_context_physRd <= lines_5_ways_0_context_physRd;
      lines_4_ways_0_context_robId <= lines_5_ways_0_context_robId;
      lines_4_ways_0_context_euCtx_0 <= lines_5_ways_0_context_euCtx_0;
      lines_4_ways_0_context_euCtx_1 <= lines_5_ways_0_context_euCtx_1;
      lines_4_ways_0_triggers <= (lines_5_ways_0_triggers >>> 1'd1);
      lines_4_ways_0_sel <= lines_5_ways_0_selComb;
      lines_5_ways_0_context_staticWake <= lines_6_ways_0_context_staticWake;
      lines_5_ways_0_context_physRd <= lines_6_ways_0_context_physRd;
      lines_5_ways_0_context_robId <= lines_6_ways_0_context_robId;
      lines_5_ways_0_context_euCtx_0 <= lines_6_ways_0_context_euCtx_0;
      lines_5_ways_0_context_euCtx_1 <= lines_6_ways_0_context_euCtx_1;
      lines_5_ways_0_triggers <= (lines_6_ways_0_triggers >>> 1'd1);
      lines_5_ways_0_sel <= lines_6_ways_0_selComb;
      lines_6_ways_0_context_staticWake <= lines_7_ways_0_context_staticWake;
      lines_6_ways_0_context_physRd <= lines_7_ways_0_context_physRd;
      lines_6_ways_0_context_robId <= lines_7_ways_0_context_robId;
      lines_6_ways_0_context_euCtx_0 <= lines_7_ways_0_context_euCtx_0;
      lines_6_ways_0_context_euCtx_1 <= lines_7_ways_0_context_euCtx_1;
      lines_6_ways_0_triggers <= (lines_7_ways_0_triggers >>> 1'd1);
      lines_6_ways_0_sel <= lines_7_ways_0_selComb;
      lines_7_ways_0_context_staticWake <= io_push_payload_slots_0_context_staticWake;
      lines_7_ways_0_context_physRd <= io_push_payload_slots_0_context_physRd;
      lines_7_ways_0_context_robId <= io_push_payload_slots_0_context_robId;
      lines_7_ways_0_context_euCtx_0 <= io_push_payload_slots_0_context_euCtx_0;
      lines_7_ways_0_context_euCtx_1 <= io_push_payload_slots_0_context_euCtx_1;
      lines_7_ways_0_triggers <= io_push_payload_slots_0_event;
      lines_7_ways_0_sel <= io_push_payload_slots_0_sel;
    end
    if(when_IssueQueue_l109) begin
      lines_0_ways_0_triggers[0] <= 1'b0;
      lines_1_ways_0_triggers[0] <= 1'b0;
      lines_2_ways_0_triggers[0] <= 1'b0;
      lines_3_ways_0_triggers[0] <= 1'b0;
      lines_4_ways_0_triggers[0] <= 1'b0;
      lines_5_ways_0_triggers[0] <= 1'b0;
      lines_6_ways_0_triggers[0] <= 1'b0;
      lines_7_ways_0_triggers[0] <= 1'b0;
    end
    if(when_IssueQueue_l109_1) begin
      lines_1_ways_0_triggers[1] <= 1'b0;
      lines_2_ways_0_triggers[1] <= 1'b0;
      lines_3_ways_0_triggers[1] <= 1'b0;
      lines_4_ways_0_triggers[1] <= 1'b0;
      lines_5_ways_0_triggers[1] <= 1'b0;
      lines_6_ways_0_triggers[1] <= 1'b0;
      lines_7_ways_0_triggers[1] <= 1'b0;
    end
    if(when_IssueQueue_l109_2) begin
      lines_2_ways_0_triggers[2] <= 1'b0;
      lines_3_ways_0_triggers[2] <= 1'b0;
      lines_4_ways_0_triggers[2] <= 1'b0;
      lines_5_ways_0_triggers[2] <= 1'b0;
      lines_6_ways_0_triggers[2] <= 1'b0;
      lines_7_ways_0_triggers[2] <= 1'b0;
    end
    if(when_IssueQueue_l109_3) begin
      lines_3_ways_0_triggers[3] <= 1'b0;
      lines_4_ways_0_triggers[3] <= 1'b0;
      lines_5_ways_0_triggers[3] <= 1'b0;
      lines_6_ways_0_triggers[3] <= 1'b0;
      lines_7_ways_0_triggers[3] <= 1'b0;
    end
    if(when_IssueQueue_l109_4) begin
      lines_4_ways_0_triggers[4] <= 1'b0;
      lines_5_ways_0_triggers[4] <= 1'b0;
      lines_6_ways_0_triggers[4] <= 1'b0;
      lines_7_ways_0_triggers[4] <= 1'b0;
    end
    if(when_IssueQueue_l109_5) begin
      lines_5_ways_0_triggers[5] <= 1'b0;
      lines_6_ways_0_triggers[5] <= 1'b0;
      lines_7_ways_0_triggers[5] <= 1'b0;
    end
    if(when_IssueQueue_l109_6) begin
      lines_6_ways_0_triggers[6] <= 1'b0;
      lines_7_ways_0_triggers[6] <= 1'b0;
    end
    if(when_IssueQueue_l109_7) begin
      lines_7_ways_0_triggers[7] <= 1'b0;
    end
    if(clear) begin
      lines_0_ways_0_sel <= 2'b00;
      lines_1_ways_0_sel <= 2'b00;
      lines_2_ways_0_sel <= 2'b00;
      lines_3_ways_0_sel <= 2'b00;
      lines_4_ways_0_sel <= 2'b00;
      lines_5_ways_0_sel <= 2'b00;
      lines_6_ways_0_sel <= 2'b00;
      lines_7_ways_0_sel <= 2'b00;
    end
  end


endmodule

module PrefetchPredictor (
  input  wire          io_learn_valid,
  input  wire [31:0]   io_learn_payload_physical,
  input  wire          io_learn_payload_allocate,
  output wire          io_prediction_cmd_valid,
  input  wire          io_prediction_cmd_ready,
  output wire [31:0]   io_prediction_cmd_payload,
  input  wire          io_prediction_rsp_valid,
  input  wire          io_prediction_rsp_payload
);


  assign io_prediction_cmd_valid = 1'b0;
  assign io_prediction_cmd_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;

endmodule

module DivRadix4 (
  input  wire          io_flush,
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [31:0]   io_cmd_payload_a,
  input  wire [31:0]   io_cmd_payload_b,
  output wire          io_rsp_valid,
  input  wire          io_rsp_ready,
  output wire [34:0]   io_rsp_payload_result,
  output wire [32:0]   io_rsp_payload_remain,
  input  wire          clk,
  input  wire          reset
);

  wire       [33:0]   _zz_div3;
  wire       [32:0]   _zz_div3_1;
  wire       [32:0]   _zz_div3_2;
  wire       [7:0]    _zz_shifter_1;
  wire       [15:0]   _zz_shifter_2;
  wire       [23:0]   _zz_shifter_3;
  reg        [3:0]    counter;
  reg                 busy;
  wire                io_rsp_fire;
  reg                 done;
  wire                when_DivRadix4_l32;
  reg        [31:0]   shifter;
  reg        [31:0]   numerator;
  reg        [31:0]   result;
  reg        [33:0]   div1;
  reg        [33:0]   div3;
  wire       [33:0]   div2;
  wire       [33:0]   shifted;
  wire       [34:0]   sub1;
  wire       [34:0]   sub2;
  wire       [34:0]   sub3;
  wire                when_DivRadix4_l51;
  reg        [33:0]   _zz_shifter;
  wire                when_DivRadix4_l55;
  wire                when_DivRadix4_l59;
  wire                when_DivRadix4_l63;
  wire                slicesZero_0;
  wire                slicesZero_1;
  wire                slicesZero_2;
  wire       [2:0]    shiftSel;
  wire       [3:0]    _zz_sel;
  wire                _zz_sel_1;
  wire                _zz_sel_2;
  wire                _zz_sel_3;
  reg        [3:0]    _zz_sel_4;
  wire       [3:0]    _zz_sel_5;
  wire                _zz_sel_6;
  wire                _zz_sel_7;
  wire                _zz_sel_8;
  wire       [1:0]    sel;
  wire                when_DivRadix4_l77;

  assign _zz_div3_1 = {1'b0,io_cmd_payload_b};
  assign _zz_div3 = {1'd0, _zz_div3_1};
  assign _zz_div3_2 = ({1'd0,io_cmd_payload_b} <<< 1'd1);
  assign _zz_shifter_1 = io_cmd_payload_a[31 : 24];
  assign _zz_shifter_2 = io_cmd_payload_a[31 : 16];
  assign _zz_shifter_3 = io_cmd_payload_a[31 : 8];
  assign io_rsp_fire = (io_rsp_valid && io_rsp_ready);
  assign when_DivRadix4_l32 = (busy && (counter == 4'b1111));
  assign div2 = (div1 <<< 1);
  assign shifted = {shifter,numerator[31 : 30]};
  assign sub1 = ({1'b0,shifted} - {1'b0,div1});
  assign sub2 = ({1'b0,shifted} - {1'b0,div2});
  assign sub3 = ({1'b0,shifted} - {1'b0,div3});
  assign io_rsp_valid = done;
  assign io_rsp_payload_result = {3'd0, result};
  assign io_rsp_payload_remain = {1'd0, shifter};
  assign io_cmd_ready = (! busy);
  assign when_DivRadix4_l51 = (! done);
  always @(*) begin
    _zz_shifter = shifted;
    if(when_DivRadix4_l55) begin
      _zz_shifter = sub1[33:0];
    end
    if(when_DivRadix4_l59) begin
      _zz_shifter = sub2[33:0];
    end
    if(when_DivRadix4_l63) begin
      _zz_shifter = sub3[33:0];
    end
  end

  assign when_DivRadix4_l55 = (! sub1[34]);
  assign when_DivRadix4_l59 = (! sub2[34]);
  assign when_DivRadix4_l63 = (! sub3[34]);
  assign slicesZero_0 = (io_cmd_payload_a[15 : 8] == 8'h00);
  assign slicesZero_1 = (io_cmd_payload_a[23 : 16] == 8'h00);
  assign slicesZero_2 = (io_cmd_payload_a[31 : 24] == 8'h00);
  assign shiftSel = {(&slicesZero_2),{(&{slicesZero_2,slicesZero_1}),(&{slicesZero_2,{slicesZero_1,slicesZero_0}})}};
  assign _zz_sel = {1'b1,shiftSel};
  assign _zz_sel_1 = _zz_sel[0];
  assign _zz_sel_2 = _zz_sel[1];
  assign _zz_sel_3 = _zz_sel[2];
  always @(*) begin
    _zz_sel_4[0] = (_zz_sel_1 && (! 1'b0));
    _zz_sel_4[1] = (_zz_sel_2 && (! _zz_sel_1));
    _zz_sel_4[2] = (_zz_sel_3 && (! (|{_zz_sel_2,_zz_sel_1})));
    _zz_sel_4[3] = (_zz_sel[3] && (! (|{_zz_sel_3,{_zz_sel_2,_zz_sel_1}})));
  end

  assign _zz_sel_5 = _zz_sel_4;
  assign _zz_sel_6 = _zz_sel_5[3];
  assign _zz_sel_7 = (_zz_sel_5[1] || _zz_sel_6);
  assign _zz_sel_8 = (_zz_sel_5[2] || _zz_sel_6);
  assign sel = {_zz_sel_8,_zz_sel_7};
  assign when_DivRadix4_l77 = (! busy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      busy <= 1'b0;
      done <= 1'b0;
    end else begin
      if(io_rsp_fire) begin
        busy <= 1'b0;
      end
      if(when_DivRadix4_l32) begin
        done <= 1'b1;
      end
      if(io_rsp_fire) begin
        done <= 1'b0;
      end
      if(when_DivRadix4_l77) begin
        busy <= io_cmd_valid;
      end
      if(io_flush) begin
        done <= 1'b0;
        busy <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(when_DivRadix4_l51) begin
      counter <= (counter + 4'b0001);
      result <= (result <<< 2);
      if(when_DivRadix4_l55) begin
        result[1 : 0] <= 2'b01;
      end
      if(when_DivRadix4_l59) begin
        result[1 : 0] <= 2'b10;
      end
      if(when_DivRadix4_l63) begin
        result[1 : 0] <= 2'b11;
      end
      shifter <= _zz_shifter[31:0];
      numerator <= (numerator <<< 2);
    end
    if(when_DivRadix4_l77) begin
      div1 <= {2'd0, io_cmd_payload_b};
      div3 <= (_zz_div3 + {1'b0,_zz_div3_2});
      result <= ((io_cmd_payload_b == 32'h00000000) ? 32'hffffffff : 32'h00000000);
      case(sel)
        2'b11 : begin
          counter <= 4'b0000;
          shifter <= 32'h00000000;
          numerator <= (io_cmd_payload_a <<< 0);
        end
        2'b10 : begin
          counter <= 4'b0100;
          shifter <= {24'd0, _zz_shifter_1};
          numerator <= (io_cmd_payload_a <<< 8);
        end
        2'b01 : begin
          counter <= 4'b1000;
          shifter <= {16'd0, _zz_shifter_2};
          numerator <= (io_cmd_payload_a <<< 16);
        end
        default : begin
          counter <= 4'b1100;
          shifter <= {8'd0, _zz_shifter_3};
          numerator <= (io_cmd_payload_a <<< 24);
        end
      endcase
    end
  end


endmodule

module StreamFifoLowLatency (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [3:0]    io_push_payload_robId,
  input  wire [0:0]    io_push_payload_mask,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [3:0]    io_pop_payload_robId,
  output wire [0:0]    io_pop_payload_mask,
  input  wire          io_flush,
  output wire [4:0]    io_occupancy,
  output wire [4:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire                fifo_io_push_ready;
  wire                fifo_io_pop_valid;
  wire       [3:0]    fifo_io_pop_payload_robId;
  wire       [0:0]    fifo_io_pop_payload_mask;
  wire       [4:0]    fifo_io_occupancy;
  wire       [4:0]    fifo_io_availability;

  StreamFifo fifo (
    .io_push_valid         (io_push_valid                 ), //i
    .io_push_ready         (fifo_io_push_ready            ), //o
    .io_push_payload_robId (io_push_payload_robId[3:0]    ), //i
    .io_push_payload_mask  (io_push_payload_mask          ), //i
    .io_pop_valid          (fifo_io_pop_valid             ), //o
    .io_pop_ready          (io_pop_ready                  ), //i
    .io_pop_payload_robId  (fifo_io_pop_payload_robId[3:0]), //o
    .io_pop_payload_mask   (fifo_io_pop_payload_mask      ), //o
    .io_flush              (io_flush                      ), //i
    .io_occupancy          (fifo_io_occupancy[4:0]        ), //o
    .io_availability       (fifo_io_availability[4:0]     ), //o
    .clk                   (clk                           ), //i
    .reset                 (reset                         )  //i
  );
  assign io_push_ready = fifo_io_push_ready;
  assign io_pop_valid = fifo_io_pop_valid;
  assign io_pop_payload_robId = fifo_io_pop_payload_robId;
  assign io_pop_payload_mask = fifo_io_pop_payload_mask;
  assign io_occupancy = fifo_io_occupancy;
  assign io_availability = fifo_io_availability;

endmodule

module DataCache (
  input  wire          io_lock_valid,
  input  wire [31:0]   io_lock_address,
  input  wire          io_load_cmd_valid,
  output wire          io_load_cmd_ready,
  input  wire [31:0]   io_load_cmd_payload_virtual,
  input  wire [1:0]    io_load_cmd_payload_size,
  input  wire          io_load_cmd_payload_redoOnDataHazard,
  input  wire          io_load_cmd_payload_unlocked,
  input  wire          io_load_cmd_payload_unique,
  input  wire [31:0]   io_load_translated_physical,
  input  wire          io_load_translated_abord,
  input  wire [2:0]    io_load_cancels,
  output wire          io_load_rsp_valid,
  output wire [31:0]   io_load_rsp_payload_data,
  output wire          io_load_rsp_payload_fault,
  output wire          io_load_rsp_payload_redo,
  output wire [1:0]    io_load_rsp_payload_refillSlot,
  output wire          io_load_rsp_payload_refillSlotAny,
  input  wire          io_store_cmd_valid,
  output wire          io_store_cmd_ready,
  input  wire [31:0]   io_store_cmd_payload_address,
  input  wire [31:0]   io_store_cmd_payload_data,
  input  wire [3:0]    io_store_cmd_payload_mask,
  input  wire          io_store_cmd_payload_generation,
  input  wire          io_store_cmd_payload_io,
  input  wire          io_store_cmd_payload_flush,
  input  wire          io_store_cmd_payload_flushFree,
  input  wire          io_store_cmd_payload_prefetch,
  output wire          io_store_rsp_valid,
  output wire          io_store_rsp_payload_fault,
  output wire          io_store_rsp_payload_redo,
  output wire [1:0]    io_store_rsp_payload_refillSlot,
  output wire          io_store_rsp_payload_refillSlotAny,
  output wire          io_store_rsp_payload_generationKo,
  output wire          io_store_rsp_payload_flush,
  output wire          io_store_rsp_payload_prefetch,
  output wire [31:0]   io_store_rsp_payload_address,
  output wire          io_store_rsp_payload_io,
  output wire          io_mem_read_cmd_valid,
  input  wire          io_mem_read_cmd_ready,
  output wire [0:0]    io_mem_read_cmd_payload_id,
  output wire [31:0]   io_mem_read_cmd_payload_address,
  input  wire          io_mem_read_rsp_valid,
  output wire          io_mem_read_rsp_ready,
  input  wire [0:0]    io_mem_read_rsp_payload_id,
  input  wire [31:0]   io_mem_read_rsp_payload_data,
  input  wire          io_mem_read_rsp_payload_error,
  output wire          io_mem_write_cmd_valid,
  input  wire          io_mem_write_cmd_ready,
  output wire          io_mem_write_cmd_payload_last,
  output wire [31:0]   io_mem_write_cmd_payload_fragment_address,
  output wire [31:0]   io_mem_write_cmd_payload_fragment_data,
  output wire [0:0]    io_mem_write_cmd_payload_fragment_id,
  input  wire          io_mem_write_rsp_valid,
  input  wire          io_mem_write_rsp_payload_error,
  input  wire [0:0]    io_mem_write_rsp_payload_id,
  output reg  [1:0]    io_refillCompletions,
  output wire          io_refillEvent,
  output wire          io_writebackEvent,
  output wire          io_writebackBusy,
  output wire          io_tagEvent,
  input  wire          clk,
  input  wire          reset
);

  reg        [31:0]   banks_0_mem_spinal_port1;
  wire       [25:0]   ways_0_mem_spinal_port1;
  wire       [25:0]   ways_0_mem_spinal_port2;
  wire       [0:0]    status_mem_spinal_port1;
  wire       [0:0]    status_mem_spinal_port2;
  reg        [31:0]   writeback_victimBuffer_spinal_port1;
  wire       [25:0]   _zz_ways_0_mem_port;
  wire                _zz_ways_0_mem_port_1;
  wire       [0:0]    _zz_status_mem_port;
  wire       [0:0]    _zz_status_loadRead_rsp_0_dirty;
  wire       [0:0]    _zz_status_storeRead_rsp_0_dirty;
  wire       [1:0]    _zz_refill_free_1;
  wire       [1:0]    _zz_refill_free_2;
  reg        [25:0]   _zz_refill_read_cmdAddress;
  reg        [31:0]   _zz_refill_read_rspAddress;
  wire       [1:0]    _zz_writeback_free_1;
  wire       [1:0]    _zz_writeback_free_2;
  reg        [31:0]   _zz_writeback_read_address;
  wire       [3:0]    _zz_writeback_read_wordIndex;
  wire       [0:0]    _zz_writeback_read_wordIndex_1;
  wire       [4:0]    _zz_writeback_victimBuffer_port;
  reg        [31:0]   _zz_writeback_write_bufferRead_payload_address;
  wire       [3:0]    _zz_writeback_write_wordIndex;
  wire       [0:0]    _zz_writeback_write_wordIndex_1;
  wire       [0:0]    _zz_when;
  wire       [0:0]    _zz_when_1;
  wire                store_pipeline_stages_0_isThrown;
  wire                store_pipeline_stages_1_isThrown;
  wire                store_pipeline_stages_2_isThrown;
  reg                 store_pipeline_stages_1_FLUSH_FREE;
  reg        [3:0]    store_pipeline_stages_1_CPU_MASK;
  reg        [31:0]   store_pipeline_stages_1_CPU_WORD;
  reg                 store_pipeline_stages_1_IO;
  reg                 store_pipeline_stages_1_FLUSH;
  reg                 store_pipeline_stages_1_PREFETCH;
  reg                 store_pipeline_stages_1_GENERATION;
  reg                 store_pipeline_stages_2_FLUSH_FREE;
  reg        [3:0]    store_pipeline_stages_2_CPU_MASK;
  reg        [31:0]   store_pipeline_stages_2_CPU_WORD;
  reg                 store_pipeline_stages_2_IO;
  wire       [1:0]    store_pipeline_stages_2_REFILL_SLOT;
  wire                store_pipeline_stages_2_REFILL_SLOT_FULL;
  reg                 store_pipeline_stages_2_WAYS_HIT;
  reg                 store_pipeline_stages_2_MISS;
  reg                 store_pipeline_stages_2_REDO;
  reg                 store_pipeline_stages_2_FLUSH;
  wire       [0:0]    store_pipeline_stages_2_WAYS_HAZARD_resulting;
  reg        [0:0]    store_pipeline_stages_2_WAYS_HITS;
  reg                 store_pipeline_stages_2_STATUS_0_dirty;
  reg                 store_pipeline_stages_2_WAYS_TAGS_0_loaded;
  reg        [23:0]   store_pipeline_stages_2_WAYS_TAGS_0_address;
  reg                 store_pipeline_stages_2_WAYS_TAGS_0_fault;
  reg                 store_pipeline_stages_2_PREFETCH;
  reg                 store_pipeline_stages_2_GENERATION;
  wire                store_pipeline_stages_2_GENERATION_OK;
  wire                store_pipeline_stages_2_PROBE;
  reg        [1:0]    store_pipeline_stages_2_REFILL_HITS_EARLY;
  wire       [1:0]    store_pipeline_stages_2_REFILL_HITS;
  reg        [1:0]    store_pipeline_stages_1_REFILL_HITS_EARLY;
  wire                store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  wire                store_pipeline_stages_1_STATUS_0_dirty;
  wire                store_pipeline_stages_1_WAYS_HIT;
  wire       [0:0]    store_pipeline_stages_1_WAYS_HITS;
  wire                store_pipeline_stages_1_WAYS_TAGS_0_loaded;
  wire       [23:0]   store_pipeline_stages_1_WAYS_TAGS_0_address;
  wire                store_pipeline_stages_1_WAYS_TAGS_0_fault;
  wire                store_pipeline_stages_1_ready;
  wire       [0:0]    store_pipeline_stages_0_WAYS_HAZARD;
  wire                store_pipeline_stages_0_GENERATION;
  wire                store_pipeline_stages_0_PREFETCH;
  wire                store_pipeline_stages_0_FLUSH_FREE;
  wire                store_pipeline_stages_0_FLUSH;
  wire                store_pipeline_stages_0_IO;
  wire       [3:0]    store_pipeline_stages_0_CPU_MASK;
  wire       [31:0]   store_pipeline_stages_0_CPU_WORD;
  wire       [31:0]   store_pipeline_stages_0_ADDRESS_POST_TRANSLATION;
  reg        [31:0]   store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  reg        [0:0]    store_pipeline_stages_2_WAYS_HAZARD;
  wire       [0:0]    store_pipeline_stages_2_WAYS_HAZARD_overloaded;
  reg        [31:0]   store_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
  reg        [0:0]    store_pipeline_stages_1_WAYS_HAZARD;
  wire       [0:0]    store_pipeline_stages_1_WAYS_HAZARD_overloaded;
  wire                load_pipeline_stages_0_isThrown;
  wire                load_pipeline_stages_1_isThrown;
  wire                load_pipeline_stages_2_isThrown;
  reg                 load_pipeline_stages_1_NEED_UNIQUE;
  wire       [1:0]    load_pipeline_stages_2_REFILL_SLOT;
  wire                load_pipeline_stages_2_REFILL_SLOT_FULL;
  reg                 load_pipeline_stages_2_ABORD;
  wire                load_pipeline_stages_2_FAULT;
  reg                 load_pipeline_stages_2_MISS;
  reg                 load_pipeline_stages_2_LOCKED;
  reg                 load_pipeline_stages_2_REDO;
  reg                 load_pipeline_stages_2_NEED_UNIQUE;
  wire       [0:0]    load_pipeline_stages_2_WAYS_HAZARD_resulting;
  reg        [0:0]    load_pipeline_stages_2_BANK_BUSY_REMAPPED;
  reg                 load_pipeline_stages_2_STATUS_0_dirty;
  reg                 load_pipeline_stages_2_WAYS_TAGS_0_loaded;
  reg        [23:0]   load_pipeline_stages_2_WAYS_TAGS_0_address;
  reg                 load_pipeline_stages_2_WAYS_TAGS_0_fault;
  reg                 load_pipeline_stages_1_UNLOCKED;
  wire                load_pipeline_stages_1_LOCKED;
  reg        [31:0]   load_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  wire       [1:0]    load_pipeline_stages_2_REFILL_HITS;
  wire                load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  wire                load_pipeline_stages_1_STATUS_0_dirty;
  wire                load_pipeline_stages_2_WAYS_HIT;
  wire       [0:0]    load_pipeline_stages_1_WAYS_HITS;
  wire                load_pipeline_stages_1_WAYS_TAGS_0_loaded;
  wire       [23:0]   load_pipeline_stages_1_WAYS_TAGS_0_address;
  wire                load_pipeline_stages_1_WAYS_TAGS_0_fault;
  wire                load_pipeline_stages_1_ready;
  wire                load_pipeline_stages_1_ABORD;
  wire       [31:0]   load_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
  reg        [31:0]   load_pipeline_stages_2_BANKS_MUXES_0;
  reg        [0:0]    load_pipeline_stages_2_WAYS_HITS;
  wire       [31:0]   load_pipeline_stages_2_CPU_WORD;
  wire       [31:0]   load_pipeline_stages_1_BANKS_MUXES_0;
  reg        [0:0]    load_pipeline_stages_1_BANK_BUSY;
  wire       [0:0]    load_pipeline_stages_1_BANK_BUSY_REMAPPED;
  wire       [31:0]   load_pipeline_stages_1_BANKS_WORDS_0;
  wire       [0:0]    load_pipeline_stages_0_BANK_BUSY_overloaded;
  wire                load_pipeline_stages_0_ready;
  wire       [0:0]    load_pipeline_stages_0_BANK_BUSY;
  wire                load_pipeline_stages_0_NEED_UNIQUE;
  wire                load_pipeline_stages_0_UNLOCKED;
  wire       [0:0]    load_pipeline_stages_0_WAYS_HAZARD;
  wire                load_pipeline_stages_0_REDO_ON_DATA_HAZARD;
  wire       [31:0]   load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION;
  reg        [31:0]   load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION;
  reg        [0:0]    load_pipeline_stages_2_WAYS_HAZARD;
  wire       [0:0]    load_pipeline_stages_2_WAYS_HAZARD_overloaded;
  reg        [31:0]   load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION;
  reg        [0:0]    load_pipeline_stages_1_WAYS_HAZARD;
  wire       [0:0]    load_pipeline_stages_1_WAYS_HAZARD_overloaded;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 banks_0_write_valid;
  reg        [5:0]    banks_0_write_payload_address;
  reg        [31:0]   banks_0_write_payload_data;
  reg        [3:0]    banks_0_write_payload_mask;
  reg                 banks_0_read_usedByWriteBack;
  reg                 banks_0_read_cmd_valid;
  reg        [5:0]    banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [31:0]   banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [0:0]    waysWrite_mask;
  reg        [1:0]    waysWrite_address;
  reg                 waysWrite_tag_loaded;
  reg        [23:0]   waysWrite_tag_address;
  reg                 waysWrite_tag_fault;
  reg        [0:0]    waysWrite_maskLast;
  reg        [1:0]    waysWrite_addressLast;
  wire                ways_0_loadRead_cmd_valid;
  wire       [1:0]    ways_0_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_0_loadRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [23:0]   ways_0_loadRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_0_loadRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [25:0]   _zz_ways_0_loadRead_rsp_loaded;
  wire                ways_0_storeRead_cmd_valid;
  wire       [1:0]    ways_0_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_0_storeRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [23:0]   ways_0_storeRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_0_storeRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [25:0]   _zz_ways_0_storeRead_rsp_loaded;
  reg                 status_write_valid;
  reg        [1:0]    status_write_payload_address;
  reg                 status_write_payload_data_0_dirty;
  wire                status_loadRead_cmd_valid;
  wire       [1:0]    status_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                status_loadRead_rsp_0_dirty /* synthesis syn_keep = 1 */ ;
  wire                status_storeRead_cmd_valid;
  wire       [1:0]    status_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                status_storeRead_rsp_0_dirty /* synthesis syn_keep = 1 */ ;
  reg                 status_writeLast_valid;
  reg        [1:0]    status_writeLast_payload_address;
  reg                 status_writeLast_payload_data_0_dirty;
  wire                wayRandom_willIncrement;
  wire                wayRandom_willClear;
  wire                wayRandom_willOverflowIfInc;
  wire                wayRandom_willOverflow;
  reg                 plru_write_valid;
  reg        [1:0]    plru_write_payload_address;
  reg                 plru_fromLoad_valid;
  wire       [1:0]    plru_fromLoad_payload_address;
  reg                 plru_fromStore_valid;
  wire       [1:0]    plru_fromStore_payload_address;
  reg        [2:0]    invalidate_counter;
  wire                invalidate_done;
  wire                invalidate_reservation_win;
  reg                 invalidate_reservation_take;
  wire                when_DataCache_l888;
  reg                 invalidate_firstEver;
  wire                when_DataCache_l897;
  reg                 refill_slots_0_valid;
  reg        [31:0]   refill_slots_0_address;
  reg                 refill_slots_0_cmdSent;
  reg        [0:0]    refill_slots_0_priority;
  reg                 refill_slots_0_loaded;
  reg        [0:0]    refill_slots_0_loadedCounter;
  wire                refill_slots_0_loadedDone;
  wire                when_DataCache_l934;
  wire                refill_slots_0_free;
  reg        [1:0]    refill_slots_0_victim;
  reg        [1:0]    refill_slots_0_writebackHazards;
  reg                 refill_slots_1_valid;
  reg        [31:0]   refill_slots_1_address;
  reg                 refill_slots_1_cmdSent;
  reg        [0:0]    refill_slots_1_priority;
  reg                 refill_slots_1_loaded;
  reg        [0:0]    refill_slots_1_loadedCounter;
  wire                refill_slots_1_loadedDone;
  wire                when_DataCache_l934_1;
  wire                refill_slots_1_free;
  reg        [1:0]    refill_slots_1_victim;
  reg        [1:0]    refill_slots_1_writebackHazards;
  wire       [1:0]    _zz_refill_free;
  wire       [1:0]    refill_free;
  wire                refill_full;
  reg                 refill_push_valid;
  reg        [31:0]   refill_push_payload_address;
  reg        [1:0]    refill_push_payload_victim;
  reg                 refill_push_payload_unique;
  reg                 refill_push_payload_data;
  reg        [31:0]   refill_pushCounter;
  wire                when_DataCache_l961;
  wire                _zz_11;
  wire                _zz_12;
  wire                when_DataCache_l961_1;
  wire                refill_read_arbiter_slotsWithId_0_0;
  wire                refill_read_arbiter_slotsWithId_1_0;
  wire       [1:0]    refill_read_arbiter_hits;
  wire                refill_read_arbiter_hit;
  reg        [1:0]    refill_read_arbiter_oh;
  wire                _zz_refill_read_arbiter_sel;
  wire       [0:0]    refill_read_arbiter_sel;
  reg        [1:0]    refill_read_arbiter_lock;
  wire                when_DataCache_l911;
  reg        [1:0]    refill_read_writebackHazards;
  wire                refill_read_writebackHazard;
  wire                io_mem_read_cmd_fire;
  wire                when_DataCache_l986;
  wire       [31:0]   refill_read_cmdAddress;
  wire                when_DataCache_l998;
  wire                when_DataCache_l998_1;
  wire       [31:0]   refill_read_rspAddress;
  (* keep , syn_keep *) reg        [3:0]    refill_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                refill_read_rspWithData;
  reg        [0:0]    refill_read_bankWriteNotif;
  reg                 refill_read_hadError;
  wire                when_DataCache_l1026;
  reg                 refill_read_fire;
  wire                refill_read_reservation_win;
  reg                 refill_read_reservation_take;
  wire                refill_read_faulty;
  wire                when_DataCache_l1037;
  reg                 writeback_slots_0_fire;
  reg                 writeback_slots_0_valid;
  reg        [31:0]   writeback_slots_0_address;
  reg        [0:0]    writeback_slots_0_priority;
  reg                 writeback_slots_0_readCmdDone;
  reg                 writeback_slots_0_victimBufferReady;
  reg                 writeback_slots_0_readRspDone;
  reg                 writeback_slots_0_writeCmdDone;
  wire                writeback_slots_0_free;
  reg                 writeback_slots_1_fire;
  reg                 writeback_slots_1_valid;
  reg        [31:0]   writeback_slots_1_address;
  reg        [0:0]    writeback_slots_1_priority;
  reg                 writeback_slots_1_readCmdDone;
  reg                 writeback_slots_1_victimBufferReady;
  reg                 writeback_slots_1_readRspDone;
  reg                 writeback_slots_1_writeCmdDone;
  wire                writeback_slots_1_free;
  wire       [1:0]    _zz_writeback_free;
  wire       [1:0]    writeback_free;
  wire                writeback_full;
  reg                 writeback_push_valid;
  reg        [31:0]   writeback_push_payload_address;
  wire                when_DataCache_l1128;
  wire                when_DataCache_l1128_1;
  wire                writeback_read_arbiter_slotsWithId_0_0;
  wire                writeback_read_arbiter_slotsWithId_1_0;
  wire       [1:0]    writeback_read_arbiter_hits;
  wire                writeback_read_arbiter_hit;
  reg        [1:0]    writeback_read_arbiter_oh;
  wire                _zz_writeback_read_arbiter_sel;
  wire       [0:0]    writeback_read_arbiter_sel;
  reg        [1:0]    writeback_read_arbiter_lock;
  wire                when_DataCache_l911_1;
  wire       [31:0]   writeback_read_address;
  (* keep , syn_keep *) reg        [3:0]    writeback_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                writeback_read_slotRead_valid;
  wire       [0:0]    writeback_read_slotRead_payload_id;
  wire                writeback_read_slotRead_payload_last;
  wire       [3:0]    writeback_read_slotRead_payload_wordIndex;
  wire                when_DataCache_l1175;
  wire                when_DataCache_l1185;
  reg                 writeback_read_slotReadLast_valid;
  reg        [0:0]    writeback_read_slotReadLast_payload_id;
  reg                 writeback_read_slotReadLast_payload_last;
  reg        [3:0]    writeback_read_slotReadLast_payload_wordIndex;
  wire       [31:0]   writeback_read_readedData;
  wire                writeback_write_arbiter_slotsWithId_0_0;
  wire                writeback_write_arbiter_slotsWithId_1_0;
  wire       [1:0]    writeback_write_arbiter_hits;
  wire                writeback_write_arbiter_hit;
  reg        [1:0]    writeback_write_arbiter_oh;
  wire                _zz_writeback_write_arbiter_sel;
  wire       [0:0]    writeback_write_arbiter_sel;
  reg        [1:0]    writeback_write_arbiter_lock;
  wire                when_DataCache_l911_2;
  (* keep , syn_keep *) reg        [3:0]    writeback_write_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                writeback_write_last;
  wire                writeback_write_bufferRead_valid;
  reg                 writeback_write_bufferRead_ready;
  wire       [0:0]    writeback_write_bufferRead_payload_id;
  wire       [31:0]   writeback_write_bufferRead_payload_address;
  wire                writeback_write_bufferRead_payload_last;
  wire                writeback_write_bufferRead_fire;
  wire                when_DataCache_l1253;
  wire                writeback_write_cmd_valid;
  wire                writeback_write_cmd_ready;
  wire       [0:0]    writeback_write_cmd_payload_id;
  wire       [31:0]   writeback_write_cmd_payload_address;
  wire                writeback_write_cmd_payload_last;
  reg                 writeback_write_bufferRead_rValid;
  reg        [0:0]    writeback_write_bufferRead_rData_id;
  reg        [31:0]   writeback_write_bufferRead_rData_address;
  reg                 writeback_write_bufferRead_rData_last;
  wire                when_Stream_l369;
  wire       [4:0]    _zz_writeback_write_word;
  wire       [31:0]   writeback_write_word;
  wire                load_pipeline_stages_0_valid;
  reg                 _zz_load_pipeline_stages_1_valid;
  reg                 load_pipeline_stages_1_valid;
  reg                 _zz_load_pipeline_stages_2_valid;
  reg                 load_pipeline_stages_2_valid;
  wire                _zz_load_pipeline_stages_0_throwRequest_DataCache_l1302;
  wire                load_pipeline_stages_0_throwRequest_DataCache_l1302;
  wire                _zz_load_pipeline_stages_1_throwRequest_DataCache_l1302;
  wire                load_pipeline_stages_1_throwRequest_DataCache_l1302;
  wire                load_pipeline_stages_2_throwRequest_DataCache_l1302;
  wire                when_DataCache_l1338;
  reg                 _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  wire                when_DataCache_l860;
  wire                when_DataCache_l863;
  wire                load_ctrl_reservation_win;
  reg                 load_ctrl_reservation_take;
  wire                _zz_refill_push_payload_victim;
  wire                load_ctrl_refillWayNeedWriteback;
  wire                load_ctrl_refillHit;
  wire                load_ctrl_refillLoaded;
  wire                load_ctrl_lineBusy;
  wire                load_ctrl_bankBusy;
  wire                load_ctrl_waysHitHazard;
  wire                load_ctrl_hitUnique;
  wire                load_ctrl_uniqueMiss;
  wire                load_ctrl_canRefill;
  wire                load_ctrl_askRefill;
  reg                 load_ctrl_askUpgrade;
  wire                load_ctrl_startRefill;
  wire                load_ctrl_startUpgrade;
  wire                when_DataCache_l1472;
  wire                when_DataCache_l1513;
  wire                when_Pipeline_l272;
  wire                when_Pipeline_l272_1;
  wire                store_pipeline_stages_0_valid;
  reg                 _zz_store_pipeline_stages_1_valid;
  reg                 store_pipeline_stages_1_valid;
  reg                 _zz_store_pipeline_stages_2_valid;
  reg                 store_pipeline_stages_2_valid;
  wire                store_pipeline_discardAll;
  wire                store_pipeline_stages_0_throwRequest_DataCache_l1552;
  wire                store_pipeline_stages_1_throwRequest_DataCache_l1552;
  wire                store_pipeline_stages_2_throwRequest_DataCache_l1552;
  reg                 store_target;
  reg                 _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  wire                when_DataCache_l860_1;
  wire                when_DataCache_l863_1;
  wire                store_refillCheckEarly_refillPushHit;
  wire                store_ctrl_reservation_win;
  reg                 store_ctrl_reservation_take;
  wire                store_ctrl_replacedWayNeedWriteback;
  wire                store_ctrl_refillHit;
  wire                store_ctrl_lineBusy;
  wire                store_ctrl_waysHitHazard;
  wire                store_ctrl_wasClean;
  wire                store_ctrl_bankBusy;
  wire                store_ctrl_hitUnique;
  wire                store_ctrl_hitFault;
  wire                store_ctrl_canRefill;
  wire                store_ctrl_askRefill;
  wire                store_ctrl_askUpgrade;
  reg                 store_ctrl_startRefill;
  reg                 store_ctrl_startUpgrade;
  reg                 store_ctrl_writeCache;
  reg                 store_ctrl_setDirty;
  wire       [0:0]    store_ctrl_needFlushs;
  wire                store_ctrl_needFlushs_bools_0;
  wire       [0:0]    _zz_store_ctrl_needFlushOh;
  wire       [0:0]    store_ctrl_needFlushOh;
  wire                _zz_15;
  wire                store_ctrl_needFlush;
  wire                store_ctrl_canFlush;
  wire                store_ctrl_startFlush;
  wire                when_DataCache_l1726;
  wire                when_DataCache_l1733;
  wire                when_DataCache_l1751;
  wire                when_DataCache_l1775;
  wire                when_DataCache_l1805;
  wire                when_Pipeline_l272_2;
  wire                when_Pipeline_l272_3;
  reg [7:0] banks_0_mem_symbol0 [0:63];
  reg [7:0] banks_0_mem_symbol1 [0:63];
  reg [7:0] banks_0_mem_symbol2 [0:63];
  reg [7:0] banks_0_mem_symbol3 [0:63];
  reg [7:0] _zz_banks_0_memsymbol_read;
  reg [7:0] _zz_banks_0_memsymbol_read_1;
  reg [7:0] _zz_banks_0_memsymbol_read_2;
  reg [7:0] _zz_banks_0_memsymbol_read_3;
  (* ram_style = "distributed" *) reg [25:0] ways_0_mem [0:3];
  (* ram_style = "distributed" *) reg [0:0] status_mem [0:3];
  reg [31:0] writeback_victimBuffer [0:31];

  assign _zz_status_loadRead_rsp_0_dirty = status_mem_spinal_port1[0 : 0];
  assign _zz_status_storeRead_rsp_0_dirty = status_mem_spinal_port2[0 : 0];
  assign _zz_refill_free_1 = (_zz_refill_free & (~ _zz_refill_free_2));
  assign _zz_refill_free_2 = (_zz_refill_free - 2'b01);
  assign _zz_writeback_free_1 = (_zz_writeback_free & (~ _zz_writeback_free_2));
  assign _zz_writeback_free_2 = (_zz_writeback_free - 2'b01);
  assign _zz_writeback_read_wordIndex_1 = writeback_read_slotRead_valid;
  assign _zz_writeback_read_wordIndex = {3'd0, _zz_writeback_read_wordIndex_1};
  assign _zz_writeback_write_wordIndex_1 = (writeback_write_bufferRead_fire && 1'b1);
  assign _zz_writeback_write_wordIndex = {3'd0, _zz_writeback_write_wordIndex_1};
  assign _zz_when = 1'b1;
  assign _zz_when_1 = 1'b1;
  assign _zz_ways_0_mem_port = {waysWrite_tag_fault,{waysWrite_tag_address,waysWrite_tag_loaded}};
  assign _zz_ways_0_mem_port_1 = waysWrite_mask[0];
  assign _zz_status_mem_port = status_write_payload_data_0_dirty;
  assign _zz_writeback_victimBuffer_port = {writeback_read_slotReadLast_payload_id,writeback_read_slotReadLast_payload_wordIndex};
  always @(*) begin
    banks_0_mem_spinal_port1 = {_zz_banks_0_memsymbol_read_3, _zz_banks_0_memsymbol_read_2, _zz_banks_0_memsymbol_read_1, _zz_banks_0_memsymbol_read};
  end
  always @(posedge clk) begin
    if(banks_0_write_payload_mask[0] && banks_0_write_valid) begin
      banks_0_mem_symbol0[banks_0_write_payload_address] <= banks_0_write_payload_data[7 : 0];
    end
    if(banks_0_write_payload_mask[1] && banks_0_write_valid) begin
      banks_0_mem_symbol1[banks_0_write_payload_address] <= banks_0_write_payload_data[15 : 8];
    end
    if(banks_0_write_payload_mask[2] && banks_0_write_valid) begin
      banks_0_mem_symbol2[banks_0_write_payload_address] <= banks_0_write_payload_data[23 : 16];
    end
    if(banks_0_write_payload_mask[3] && banks_0_write_valid) begin
      banks_0_mem_symbol3[banks_0_write_payload_address] <= banks_0_write_payload_data[31 : 24];
    end
  end

  always @(posedge clk) begin
    if(banks_0_read_cmd_valid) begin
      _zz_banks_0_memsymbol_read <= banks_0_mem_symbol0[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_1 <= banks_0_mem_symbol1[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_2 <= banks_0_mem_symbol2[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_3 <= banks_0_mem_symbol3[banks_0_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_ways_0_mem_port_1) begin
      ways_0_mem[waysWrite_address] <= _zz_ways_0_mem_port;
    end
  end

  assign ways_0_mem_spinal_port1 = ways_0_mem[ways_0_loadRead_cmd_payload];
  assign ways_0_mem_spinal_port2 = ways_0_mem[ways_0_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_2) begin
      status_mem[status_write_payload_address] <= _zz_status_mem_port;
    end
  end

  assign status_mem_spinal_port1 = status_mem[status_loadRead_cmd_payload];
  assign status_mem_spinal_port2 = status_mem[status_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_1) begin
      writeback_victimBuffer[_zz_writeback_victimBuffer_port] <= writeback_read_readedData;
    end
  end

  always @(posedge clk) begin
    if(writeback_write_bufferRead_ready) begin
      writeback_victimBuffer_spinal_port1 <= writeback_victimBuffer[_zz_writeback_write_word];
    end
  end

  always @(*) begin
    case(refill_read_arbiter_sel)
      1'b0 : _zz_refill_read_cmdAddress = refill_slots_0_address[31 : 6];
      default : _zz_refill_read_cmdAddress = refill_slots_1_address[31 : 6];
    endcase
  end

  always @(*) begin
    case(io_mem_read_rsp_payload_id)
      1'b0 : _zz_refill_read_rspAddress = refill_slots_0_address;
      default : _zz_refill_read_rspAddress = refill_slots_1_address;
    endcase
  end

  always @(*) begin
    case(writeback_read_arbiter_sel)
      1'b0 : _zz_writeback_read_address = writeback_slots_0_address;
      default : _zz_writeback_read_address = writeback_slots_1_address;
    endcase
  end

  always @(*) begin
    case(writeback_write_arbiter_sel)
      1'b0 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_0_address;
      default : _zz_writeback_write_bufferRead_payload_address = writeback_slots_1_address;
    endcase
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(writeback_read_slotReadLast_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(status_write_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    banks_0_read_usedByWriteBack = 1'b0;
    if(when_DataCache_l1185) begin
      banks_0_read_usedByWriteBack = 1'b1;
    end
  end

  assign banks_0_read_rsp = banks_0_mem_spinal_port1;
  always @(*) begin
    banks_0_read_cmd_valid = 1'b0;
    if(when_DataCache_l1185) begin
      banks_0_read_cmd_valid = 1'b1;
    end
    if(when_DataCache_l1338) begin
      banks_0_read_cmd_valid = (! (load_pipeline_stages_0_valid && (! load_pipeline_stages_0_ready)));
    end
  end

  always @(*) begin
    banks_0_read_cmd_payload = 6'bxxxxxx;
    if(when_DataCache_l1185) begin
      banks_0_read_cmd_payload = {writeback_read_address[7 : 6],writeback_read_wordIndex};
    end
    if(when_DataCache_l1338) begin
      banks_0_read_cmd_payload = load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION[7 : 2];
    end
  end

  always @(*) begin
    waysWrite_mask = 1'b0;
    if(when_DataCache_l888) begin
      waysWrite_mask = 1'b1;
    end
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        waysWrite_mask[0] = 1'b1;
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_mask[0] = 1'b1;
    end
    if(when_DataCache_l1751) begin
      waysWrite_mask[0] = 1'b1;
    end
    if(store_ctrl_startFlush) begin
      if(store_pipeline_stages_2_FLUSH_FREE) begin
        if(_zz_15) begin
          waysWrite_mask[0] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    waysWrite_address = 2'bxx;
    if(when_DataCache_l888) begin
      waysWrite_address = invalidate_counter[1:0];
    end
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        waysWrite_address = refill_read_rspAddress[7 : 6];
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_address = load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[7 : 6];
    end
    if(when_DataCache_l1751) begin
      waysWrite_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 6];
    end
    if(store_ctrl_startFlush) begin
      waysWrite_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 6];
    end
  end

  always @(*) begin
    waysWrite_tag_loaded = 1'bx;
    if(when_DataCache_l888) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        waysWrite_tag_loaded = 1'b1;
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(when_DataCache_l1751) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(store_ctrl_startFlush) begin
      waysWrite_tag_loaded = 1'b0;
    end
  end

  always @(*) begin
    waysWrite_tag_address = 24'bxxxxxxxxxxxxxxxxxxxxxxxx;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        waysWrite_tag_address = refill_read_rspAddress[31 : 8];
      end
    end
  end

  always @(*) begin
    waysWrite_tag_fault = 1'bx;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        waysWrite_tag_fault = refill_read_faulty;
      end
    end
  end

  assign _zz_ways_0_loadRead_rsp_loaded = ways_0_mem_spinal_port1;
  assign ways_0_loadRead_rsp_loaded = _zz_ways_0_loadRead_rsp_loaded[0];
  assign ways_0_loadRead_rsp_address = _zz_ways_0_loadRead_rsp_loaded[24 : 1];
  assign ways_0_loadRead_rsp_fault = _zz_ways_0_loadRead_rsp_loaded[25];
  assign _zz_ways_0_storeRead_rsp_loaded = ways_0_mem_spinal_port2;
  assign ways_0_storeRead_rsp_loaded = _zz_ways_0_storeRead_rsp_loaded[0];
  assign ways_0_storeRead_rsp_address = _zz_ways_0_storeRead_rsp_loaded[24 : 1];
  assign ways_0_storeRead_rsp_fault = _zz_ways_0_storeRead_rsp_loaded[25];
  always @(*) begin
    status_write_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      status_write_valid = 1'b1;
    end
    if(when_DataCache_l1726) begin
      status_write_valid = 1'b1;
    end
  end

  always @(*) begin
    status_write_payload_address = 2'bxx;
    if(load_ctrl_startRefill) begin
      status_write_payload_address = load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[7 : 6];
    end
    if(when_DataCache_l1726) begin
      status_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 6];
    end
  end

  always @(*) begin
    status_write_payload_data_0_dirty = 1'bx;
    if(load_ctrl_startRefill) begin
      status_write_payload_data_0_dirty = load_pipeline_stages_2_STATUS_0_dirty;
      if(_zz_when[0]) begin
        status_write_payload_data_0_dirty = 1'b0;
      end
    end
    if(when_DataCache_l1726) begin
      status_write_payload_data_0_dirty = store_pipeline_stages_2_STATUS_0_dirty;
    end
    if(when_DataCache_l1751) begin
      status_write_payload_data_0_dirty = 1'b0;
    end
    if(store_ctrl_setDirty) begin
      if(store_pipeline_stages_2_WAYS_HITS[0]) begin
        status_write_payload_data_0_dirty = 1'b1;
      end
    end
    if(store_ctrl_startFlush) begin
      if(_zz_15) begin
        status_write_payload_data_0_dirty = 1'b0;
      end
    end
  end

  assign status_loadRead_rsp_0_dirty = _zz_status_loadRead_rsp_0_dirty[0];
  assign status_storeRead_rsp_0_dirty = _zz_status_storeRead_rsp_0_dirty[0];
  assign wayRandom_willClear = 1'b0;
  assign wayRandom_willOverflowIfInc = 1'b1;
  assign wayRandom_willOverflow = (wayRandom_willOverflowIfInc && wayRandom_willIncrement);
  assign wayRandom_willIncrement = 1'b1;
  always @(*) begin
    plru_write_valid = (plru_fromLoad_valid || plru_fromStore_valid);
    if(when_DataCache_l897) begin
      plru_write_valid = 1'b1;
    end
  end

  always @(*) begin
    plru_write_payload_address = (plru_fromLoad_valid ? plru_fromLoad_payload_address : plru_fromStore_payload_address);
    if(when_DataCache_l897) begin
      plru_write_payload_address = invalidate_counter[1:0];
    end
  end

  assign invalidate_done = invalidate_counter[2];
  always @(*) begin
    invalidate_reservation_take = 1'b0;
    if(when_DataCache_l888) begin
      invalidate_reservation_take = 1'b1;
    end
  end

  assign when_DataCache_l888 = ((! invalidate_done) && invalidate_reservation_win);
  assign when_DataCache_l897 = ((! invalidate_done) && invalidate_firstEver);
  assign refill_slots_0_loadedDone = (refill_slots_0_loadedCounter == 1'b1);
  assign when_DataCache_l934 = (refill_slots_0_loadedDone && 1'b1);
  assign refill_slots_0_free = (! refill_slots_0_valid);
  assign refill_slots_1_loadedDone = (refill_slots_1_loadedCounter == 1'b1);
  assign when_DataCache_l934_1 = (refill_slots_1_loadedDone && 1'b1);
  assign refill_slots_1_free = (! refill_slots_1_valid);
  assign _zz_refill_free = {refill_slots_1_free,refill_slots_0_free};
  assign refill_free = {_zz_refill_free_1[1],refill_slots_0_free};
  assign refill_full = (&{(! refill_slots_1_free),(! refill_slots_0_free)});
  always @(*) begin
    refill_push_valid = 1'b0;
    if(when_DataCache_l1472) begin
      refill_push_valid = 1'b1;
    end
    if(when_DataCache_l1751) begin
      refill_push_valid = 1'b1;
    end
  end

  always @(*) begin
    refill_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_DataCache_l1472) begin
      refill_push_payload_address = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
    end
    if(when_DataCache_l1751) begin
      refill_push_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
    end
  end

  always @(*) begin
    refill_push_payload_victim = 2'bxx;
    if(load_ctrl_askUpgrade) begin
      refill_push_payload_victim = 2'b00;
    end else begin
      refill_push_payload_victim = ((load_ctrl_refillWayNeedWriteback && _zz_refill_push_payload_victim) ? writeback_free : 2'b00);
    end
    if(when_DataCache_l1751) begin
      refill_push_payload_victim = (((store_ctrl_replacedWayNeedWriteback && store_ctrl_askRefill) && store_pipeline_stages_2_STATUS_0_dirty) ? writeback_free : 2'b00);
    end
  end

  always @(*) begin
    refill_push_payload_unique = 1'bx;
    if(when_DataCache_l1472) begin
      refill_push_payload_unique = load_pipeline_stages_2_NEED_UNIQUE;
    end
    if(when_DataCache_l1751) begin
      refill_push_payload_unique = 1'b1;
    end
  end

  always @(*) begin
    refill_push_payload_data = 1'bx;
    if(when_DataCache_l1472) begin
      refill_push_payload_data = load_ctrl_askRefill;
    end
    if(when_DataCache_l1751) begin
      refill_push_payload_data = store_ctrl_askRefill;
    end
  end

  assign when_DataCache_l961 = refill_free[0];
  assign _zz_11 = refill_free[0];
  assign _zz_12 = refill_free[1];
  assign when_DataCache_l961_1 = refill_free[1];
  assign refill_read_arbiter_slotsWithId_0_0 = (((refill_slots_0_valid && (! refill_slots_0_cmdSent)) && (refill_slots_0_victim == 2'b00)) && (refill_slots_0_writebackHazards == 2'b00));
  assign refill_read_arbiter_slotsWithId_1_0 = (((refill_slots_1_valid && (! refill_slots_1_cmdSent)) && (refill_slots_1_victim == 2'b00)) && (refill_slots_1_writebackHazards == 2'b00));
  assign refill_read_arbiter_hits = {refill_read_arbiter_slotsWithId_1_0,refill_read_arbiter_slotsWithId_0_0};
  assign refill_read_arbiter_hit = (|refill_read_arbiter_hits);
  always @(*) begin
    refill_read_arbiter_oh = (refill_read_arbiter_hits & {((refill_read_arbiter_hits[0] & refill_slots_1_priority) == 1'b0),((refill_read_arbiter_hits[1] & refill_slots_0_priority) == 1'b0)});
    if(when_DataCache_l911) begin
      refill_read_arbiter_oh = refill_read_arbiter_lock;
    end
  end

  assign _zz_refill_read_arbiter_sel = refill_read_arbiter_oh[1];
  assign refill_read_arbiter_sel = _zz_refill_read_arbiter_sel;
  assign when_DataCache_l911 = (|refill_read_arbiter_lock);
  assign refill_read_writebackHazard = (|refill_read_writebackHazards);
  assign io_mem_read_cmd_fire = (io_mem_read_cmd_valid && io_mem_read_cmd_ready);
  assign when_DataCache_l986 = (io_mem_read_cmd_fire || refill_read_writebackHazard);
  assign refill_read_cmdAddress = {_zz_refill_read_cmdAddress,6'h00};
  assign io_mem_read_cmd_valid = (refill_read_arbiter_hit && (! refill_read_writebackHazard));
  assign io_mem_read_cmd_payload_id = refill_read_arbiter_sel;
  assign io_mem_read_cmd_payload_address = refill_read_cmdAddress;
  assign when_DataCache_l998 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_DataCache_l998_1 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign refill_read_rspAddress = _zz_refill_read_rspAddress;
  assign refill_read_rspWithData = 1'b1;
  always @(*) begin
    refill_read_bankWriteNotif = 1'b0;
    refill_read_bankWriteNotif[0] = ((io_mem_read_rsp_valid && refill_read_rspWithData) && 1'b1);
  end

  always @(*) begin
    banks_0_write_valid = refill_read_bankWriteNotif[0];
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1775) begin
        banks_0_write_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_address = {refill_read_rspAddress[7 : 6],refill_read_wordIndex};
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1775) begin
        banks_0_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 2];
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_data = io_mem_read_rsp_payload_data;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1775) begin
        banks_0_write_payload_data[31 : 0] = store_pipeline_stages_2_CPU_WORD;
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_mask = 4'b1111;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1775) begin
        banks_0_write_payload_mask = 4'b0000;
        if(_zz_when_1[0]) begin
          banks_0_write_payload_mask[3 : 0] = store_pipeline_stages_2_CPU_MASK;
        end
      end
    end
  end

  assign when_DataCache_l1026 = (io_mem_read_rsp_valid && io_mem_read_rsp_payload_error);
  always @(*) begin
    refill_read_fire = 1'b0;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        refill_read_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    refill_read_reservation_take = 1'b0;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        refill_read_reservation_take = 1'b1;
      end
    end
  end

  assign refill_read_faulty = (refill_read_hadError || io_mem_read_rsp_payload_error);
  always @(*) begin
    io_refillCompletions = 2'b00;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        io_refillCompletions[io_mem_read_rsp_payload_id] = 1'b1;
      end
    end
  end

  assign io_mem_read_rsp_ready = 1'b1;
  assign when_DataCache_l1037 = ((refill_read_wordIndex == 4'b1111) || (! refill_read_rspWithData));
  always @(*) begin
    writeback_slots_0_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        1'b0 : begin
          writeback_slots_0_fire = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_0_free = (! writeback_slots_0_valid);
  always @(*) begin
    refill_read_writebackHazards[0] = (writeback_slots_0_valid && (writeback_slots_0_address[31 : 6] == refill_read_cmdAddress[31 : 6]));
    refill_read_writebackHazards[1] = (writeback_slots_1_valid && (writeback_slots_1_address[31 : 6] == refill_read_cmdAddress[31 : 6]));
  end

  always @(*) begin
    writeback_slots_1_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        1'b0 : begin
        end
        default : begin
          writeback_slots_1_fire = 1'b1;
        end
      endcase
    end
  end

  assign writeback_slots_1_free = (! writeback_slots_1_valid);
  assign io_writebackBusy = (|{writeback_slots_1_valid,writeback_slots_0_valid});
  assign _zz_writeback_free = {writeback_slots_1_free,writeback_slots_0_free};
  assign writeback_free = {_zz_writeback_free_1[1],writeback_slots_0_free};
  assign writeback_full = (&{(! writeback_slots_1_free),(! writeback_slots_0_free)});
  always @(*) begin
    writeback_push_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      writeback_push_valid = load_ctrl_refillWayNeedWriteback;
    end
    if(when_DataCache_l1733) begin
      writeback_push_valid = (store_ctrl_replacedWayNeedWriteback || store_ctrl_startFlush);
    end
  end

  always @(*) begin
    writeback_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(load_ctrl_startRefill) begin
      writeback_push_payload_address = ({6'd0,{load_pipeline_stages_2_WAYS_TAGS_0_address,load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[7 : 6]}} <<< 3'd6);
    end
    if(when_DataCache_l1733) begin
      writeback_push_payload_address = ({6'd0,{store_pipeline_stages_2_WAYS_TAGS_0_address,store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 6]}} <<< 3'd6);
    end
  end

  assign when_DataCache_l1128 = writeback_free[0];
  assign when_DataCache_l1128_1 = writeback_free[1];
  assign writeback_read_arbiter_slotsWithId_0_0 = (writeback_slots_0_valid && (! writeback_slots_0_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_1_0 = (writeback_slots_1_valid && (! writeback_slots_1_readCmdDone));
  assign writeback_read_arbiter_hits = {writeback_read_arbiter_slotsWithId_1_0,writeback_read_arbiter_slotsWithId_0_0};
  assign writeback_read_arbiter_hit = (|writeback_read_arbiter_hits);
  always @(*) begin
    writeback_read_arbiter_oh = (writeback_read_arbiter_hits & {((writeback_read_arbiter_hits[0] & writeback_slots_1_priority) == 1'b0),((writeback_read_arbiter_hits[1] & writeback_slots_0_priority) == 1'b0)});
    if(when_DataCache_l911_1) begin
      writeback_read_arbiter_oh = writeback_read_arbiter_lock;
    end
  end

  assign _zz_writeback_read_arbiter_sel = writeback_read_arbiter_oh[1];
  assign writeback_read_arbiter_sel = _zz_writeback_read_arbiter_sel;
  assign when_DataCache_l911_1 = (|writeback_read_arbiter_lock);
  assign writeback_read_address = _zz_writeback_read_address;
  assign writeback_read_slotRead_valid = writeback_read_arbiter_hit;
  assign writeback_read_slotRead_payload_id = writeback_read_arbiter_sel;
  assign writeback_read_slotRead_payload_wordIndex = writeback_read_wordIndex;
  assign writeback_read_slotRead_payload_last = (writeback_read_wordIndex == 4'b1111);
  assign when_DataCache_l1175 = (writeback_read_slotRead_valid && writeback_read_slotRead_payload_last);
  assign when_DataCache_l1185 = (writeback_read_slotRead_valid && 1'b1);
  assign writeback_read_readedData = banks_0_read_rsp;
  assign writeback_write_arbiter_slotsWithId_0_0 = ((writeback_slots_0_valid && writeback_slots_0_victimBufferReady) && (! writeback_slots_0_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_1_0 = ((writeback_slots_1_valid && writeback_slots_1_victimBufferReady) && (! writeback_slots_1_writeCmdDone));
  assign writeback_write_arbiter_hits = {writeback_write_arbiter_slotsWithId_1_0,writeback_write_arbiter_slotsWithId_0_0};
  assign writeback_write_arbiter_hit = (|writeback_write_arbiter_hits);
  always @(*) begin
    writeback_write_arbiter_oh = (writeback_write_arbiter_hits & {((writeback_write_arbiter_hits[0] & writeback_slots_1_priority) == 1'b0),((writeback_write_arbiter_hits[1] & writeback_slots_0_priority) == 1'b0)});
    if(when_DataCache_l911_2) begin
      writeback_write_arbiter_oh = writeback_write_arbiter_lock;
    end
  end

  assign _zz_writeback_write_arbiter_sel = writeback_write_arbiter_oh[1];
  assign writeback_write_arbiter_sel = _zz_writeback_write_arbiter_sel;
  assign when_DataCache_l911_2 = (|writeback_write_arbiter_lock);
  assign writeback_write_last = (writeback_write_wordIndex == 4'b1111);
  assign writeback_write_bufferRead_valid = writeback_write_arbiter_hit;
  assign writeback_write_bufferRead_payload_id = writeback_write_arbiter_sel;
  assign writeback_write_bufferRead_payload_last = writeback_write_last;
  assign writeback_write_bufferRead_payload_address = _zz_writeback_write_bufferRead_payload_address;
  assign writeback_write_bufferRead_fire = (writeback_write_bufferRead_valid && writeback_write_bufferRead_ready);
  assign when_DataCache_l1253 = (writeback_write_bufferRead_fire && writeback_write_last);
  always @(*) begin
    writeback_write_bufferRead_ready = writeback_write_cmd_ready;
    if(when_Stream_l369) begin
      writeback_write_bufferRead_ready = 1'b1;
    end
  end

  assign when_Stream_l369 = (! writeback_write_cmd_valid);
  assign writeback_write_cmd_valid = writeback_write_bufferRead_rValid;
  assign writeback_write_cmd_payload_id = writeback_write_bufferRead_rData_id;
  assign writeback_write_cmd_payload_address = writeback_write_bufferRead_rData_address;
  assign writeback_write_cmd_payload_last = writeback_write_bufferRead_rData_last;
  assign _zz_writeback_write_word = {writeback_write_bufferRead_payload_id,writeback_write_wordIndex};
  assign writeback_write_word = writeback_victimBuffer_spinal_port1;
  assign io_mem_write_cmd_valid = writeback_write_cmd_valid;
  assign writeback_write_cmd_ready = io_mem_write_cmd_ready;
  assign io_mem_write_cmd_payload_fragment_address = writeback_write_cmd_payload_address;
  assign io_mem_write_cmd_payload_fragment_data = writeback_write_word;
  assign io_mem_write_cmd_payload_fragment_id = writeback_write_cmd_payload_id;
  assign io_mem_write_cmd_payload_last = writeback_write_cmd_payload_last;
  assign _zz_load_pipeline_stages_0_throwRequest_DataCache_l1302 = io_load_cancels[0];
  assign load_pipeline_stages_0_throwRequest_DataCache_l1302 = _zz_load_pipeline_stages_0_throwRequest_DataCache_l1302;
  assign _zz_load_pipeline_stages_1_throwRequest_DataCache_l1302 = io_load_cancels[1];
  assign load_pipeline_stages_1_throwRequest_DataCache_l1302 = _zz_load_pipeline_stages_1_throwRequest_DataCache_l1302;
  assign load_pipeline_stages_2_throwRequest_DataCache_l1302 = io_load_cancels[2];
  assign load_pipeline_stages_1_WAYS_HAZARD_overloaded = (load_pipeline_stages_1_WAYS_HAZARD | ((waysWrite_addressLast == load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[7 : 6]) ? waysWrite_maskLast : 1'b0));
  assign load_pipeline_stages_2_WAYS_HAZARD_overloaded = (load_pipeline_stages_2_WAYS_HAZARD | ((waysWrite_addressLast == load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[7 : 6]) ? waysWrite_maskLast : 1'b0));
  assign io_load_cmd_ready = 1'b1;
  assign load_pipeline_stages_0_valid = io_load_cmd_valid;
  assign load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION = io_load_cmd_payload_virtual;
  assign load_pipeline_stages_0_REDO_ON_DATA_HAZARD = io_load_cmd_payload_redoOnDataHazard;
  assign load_pipeline_stages_0_WAYS_HAZARD = 1'b0;
  assign load_pipeline_stages_0_UNLOCKED = io_load_cmd_payload_unlocked;
  assign load_pipeline_stages_0_NEED_UNIQUE = io_load_cmd_payload_unique;
  assign load_pipeline_stages_0_BANK_BUSY[0] = banks_0_read_usedByWriteBack;
  assign when_DataCache_l1338 = (! load_pipeline_stages_0_BANK_BUSY[0]);
  assign load_pipeline_stages_0_BANK_BUSY_overloaded[0] = (load_pipeline_stages_0_BANK_BUSY[0] || (banks_0_write_valid && load_pipeline_stages_0_REDO_ON_DATA_HAZARD));
  assign load_pipeline_stages_1_BANKS_WORDS_0 = banks_0_read_rsp;
  assign load_pipeline_stages_1_BANK_BUSY_REMAPPED[0] = load_pipeline_stages_1_BANK_BUSY[0];
  assign load_pipeline_stages_1_BANKS_MUXES_0 = load_pipeline_stages_1_BANKS_WORDS_0[31 : 0];
  assign load_pipeline_stages_2_CPU_WORD = (load_pipeline_stages_2_WAYS_HITS[0] ? load_pipeline_stages_2_BANKS_MUXES_0 : 32'h00000000);
  assign load_pipeline_stages_1_ADDRESS_POST_TRANSLATION = io_load_translated_physical;
  assign load_pipeline_stages_1_ABORD = io_load_translated_abord;
  assign ways_0_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign ways_0_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[7 : 6];
  assign load_pipeline_stages_1_WAYS_TAGS_0_loaded = ways_0_loadRead_rsp_loaded;
  assign load_pipeline_stages_1_WAYS_TAGS_0_address = ways_0_loadRead_rsp_address;
  assign load_pipeline_stages_1_WAYS_TAGS_0_fault = ways_0_loadRead_rsp_fault;
  assign load_pipeline_stages_1_WAYS_HITS[0] = (load_pipeline_stages_1_WAYS_TAGS_0_loaded && (load_pipeline_stages_1_WAYS_TAGS_0_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 8]));
  assign load_pipeline_stages_2_WAYS_HIT = (|load_pipeline_stages_2_WAYS_HITS);
  assign status_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign status_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[7 : 6];
  assign load_pipeline_stages_1_STATUS_0_dirty = status_loadRead_rsp_0_dirty;
  always @(*) begin
    _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = load_pipeline_stages_1_STATUS_0_dirty;
    if(when_DataCache_l860) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = status_writeLast_payload_data_0_dirty;
    end
    if(when_DataCache_l863) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = status_write_payload_data_0_dirty;
    end
  end

  assign when_DataCache_l860 = (status_writeLast_valid && (status_writeLast_payload_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[7 : 6]));
  assign when_DataCache_l863 = (status_write_valid && (status_write_payload_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[7 : 6]));
  assign load_pipeline_stages_1_STATUS_overloaded_0_dirty = _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  assign load_pipeline_stages_2_REFILL_HITS = {(refill_slots_1_valid && (refill_slots_1_address[31 : 6] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[31 : 6])),(refill_slots_0_valid && (refill_slots_0_address[31 : 6] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[31 : 6]))};
  assign load_pipeline_stages_1_LOCKED = (((! load_pipeline_stages_1_UNLOCKED) && io_lock_valid) && (io_lock_address[7 : 6] == load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[7 : 6]));
  always @(*) begin
    plru_fromLoad_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      plru_fromLoad_valid = 1'b1;
    end
    if(when_DataCache_l1513) begin
      plru_fromLoad_valid = 1'b1;
    end
  end

  assign plru_fromLoad_payload_address = load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[7 : 6];
  always @(*) begin
    load_ctrl_reservation_take = 1'b0;
    if(when_DataCache_l1472) begin
      load_ctrl_reservation_take = 1'b1;
    end
  end

  assign _zz_refill_push_payload_victim = load_pipeline_stages_2_STATUS_0_dirty;
  assign load_ctrl_refillWayNeedWriteback = (load_pipeline_stages_2_WAYS_TAGS_0_loaded && _zz_refill_push_payload_victim);
  assign load_ctrl_refillHit = (|load_pipeline_stages_2_REFILL_HITS);
  assign load_ctrl_refillLoaded = (|({refill_slots_1_loaded,refill_slots_0_loaded} & load_pipeline_stages_2_REFILL_HITS));
  assign load_ctrl_lineBusy = ((|{(refill_slots_1_valid && (refill_slots_1_address[7 : 6] == load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[7 : 6])),(refill_slots_0_valid && (refill_slots_0_address[7 : 6] == load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[7 : 6]))}) || 1'b0);
  assign load_ctrl_bankBusy = ((load_pipeline_stages_2_BANK_BUSY_REMAPPED & load_pipeline_stages_2_WAYS_HITS) != 1'b0);
  assign load_ctrl_waysHitHazard = (|(load_pipeline_stages_2_WAYS_HITS & load_pipeline_stages_2_WAYS_HAZARD_resulting));
  assign load_ctrl_hitUnique = 1'b1;
  assign load_ctrl_uniqueMiss = (load_pipeline_stages_2_NEED_UNIQUE && (! load_ctrl_hitUnique));
  always @(*) begin
    load_pipeline_stages_2_REDO = ((((((! load_pipeline_stages_2_WAYS_HIT) || load_ctrl_waysHitHazard) || load_ctrl_bankBusy) || load_ctrl_refillHit) || load_pipeline_stages_2_LOCKED) || load_ctrl_uniqueMiss);
    if(load_pipeline_stages_2_ABORD) begin
      load_pipeline_stages_2_REDO = 1'b0;
    end
  end

  always @(*) begin
    load_pipeline_stages_2_MISS = ((((! load_pipeline_stages_2_WAYS_HIT) && (! load_ctrl_waysHitHazard)) && (! load_ctrl_refillHit)) && (! load_pipeline_stages_2_LOCKED));
    if(load_pipeline_stages_2_ABORD) begin
      load_pipeline_stages_2_MISS = 1'b0;
    end
  end

  assign load_pipeline_stages_2_FAULT = (|(load_pipeline_stages_2_WAYS_HITS & load_pipeline_stages_2_WAYS_TAGS_0_fault));
  assign load_ctrl_canRefill = (((((! refill_full) && (! load_ctrl_lineBusy)) && load_ctrl_reservation_win) && (! (load_ctrl_refillWayNeedWriteback && writeback_full))) && (! load_pipeline_stages_2_WAYS_HAZARD_resulting[0]));
  assign load_ctrl_askRefill = ((load_pipeline_stages_2_MISS && load_ctrl_canRefill) && (! load_ctrl_refillHit));
  always @(*) begin
    load_ctrl_askUpgrade = (((! load_pipeline_stages_2_MISS) && load_ctrl_canRefill) && load_ctrl_uniqueMiss);
    if(load_pipeline_stages_2_ABORD) begin
      load_ctrl_askUpgrade = 1'b0;
    end
  end

  assign load_ctrl_startRefill = (load_pipeline_stages_2_valid && load_ctrl_askRefill);
  assign load_ctrl_startUpgrade = (load_pipeline_stages_2_valid && load_ctrl_askUpgrade);
  assign when_DataCache_l1472 = (load_ctrl_startRefill || load_ctrl_startUpgrade);
  assign when_DataCache_l1513 = ((load_pipeline_stages_2_valid && (! load_pipeline_stages_2_REDO)) && (! load_pipeline_stages_2_MISS));
  assign load_pipeline_stages_2_REFILL_SLOT_FULL = ((load_pipeline_stages_2_MISS && (! load_ctrl_refillHit)) && refill_full);
  assign load_pipeline_stages_2_REFILL_SLOT = (((! load_ctrl_refillLoaded) ? load_pipeline_stages_2_REFILL_HITS : 2'b00) | (load_ctrl_askRefill ? refill_free : 2'b00));
  assign io_load_rsp_valid = load_pipeline_stages_2_valid;
  assign io_load_rsp_payload_data = load_pipeline_stages_2_CPU_WORD;
  assign io_load_rsp_payload_fault = load_pipeline_stages_2_FAULT;
  assign io_load_rsp_payload_redo = load_pipeline_stages_2_REDO;
  assign io_load_rsp_payload_refillSlotAny = load_pipeline_stages_2_REFILL_SLOT_FULL;
  assign io_load_rsp_payload_refillSlot = load_pipeline_stages_2_REFILL_SLOT;
  assign load_pipeline_stages_2_isThrown = load_pipeline_stages_2_throwRequest_DataCache_l1302;
  assign load_pipeline_stages_1_isThrown = load_pipeline_stages_1_throwRequest_DataCache_l1302;
  assign load_pipeline_stages_0_isThrown = load_pipeline_stages_0_throwRequest_DataCache_l1302;
  always @(*) begin
    _zz_load_pipeline_stages_1_valid = load_pipeline_stages_0_valid;
    if(when_Pipeline_l272) begin
      _zz_load_pipeline_stages_1_valid = 1'b0;
    end
  end

  assign load_pipeline_stages_0_ready = 1'b1;
  assign when_Pipeline_l272 = (|_zz_load_pipeline_stages_0_throwRequest_DataCache_l1302);
  always @(*) begin
    _zz_load_pipeline_stages_2_valid = load_pipeline_stages_1_valid;
    if(when_Pipeline_l272_1) begin
      _zz_load_pipeline_stages_2_valid = 1'b0;
    end
  end

  assign load_pipeline_stages_1_ready = 1'b1;
  assign when_Pipeline_l272_1 = (|_zz_load_pipeline_stages_1_throwRequest_DataCache_l1302);
  assign load_pipeline_stages_2_WAYS_HAZARD_resulting = load_pipeline_stages_2_WAYS_HAZARD_overloaded;
  assign store_pipeline_discardAll = 1'b0;
  assign store_pipeline_stages_0_throwRequest_DataCache_l1552 = store_pipeline_discardAll;
  assign store_pipeline_stages_1_throwRequest_DataCache_l1552 = store_pipeline_discardAll;
  assign store_pipeline_stages_2_throwRequest_DataCache_l1552 = store_pipeline_discardAll;
  assign store_pipeline_stages_1_WAYS_HAZARD_overloaded = (store_pipeline_stages_1_WAYS_HAZARD | ((waysWrite_addressLast == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[7 : 6]) ? waysWrite_maskLast : 1'b0));
  assign store_pipeline_stages_2_WAYS_HAZARD_overloaded = (store_pipeline_stages_2_WAYS_HAZARD | ((waysWrite_addressLast == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 6]) ? waysWrite_maskLast : 1'b0));
  assign store_pipeline_stages_0_valid = io_store_cmd_valid;
  assign store_pipeline_stages_0_ADDRESS_POST_TRANSLATION = io_store_cmd_payload_address;
  assign store_pipeline_stages_0_CPU_WORD = io_store_cmd_payload_data;
  assign store_pipeline_stages_0_CPU_MASK = io_store_cmd_payload_mask;
  assign store_pipeline_stages_0_IO = (io_store_cmd_payload_io && (! io_store_cmd_payload_flush));
  assign store_pipeline_stages_0_FLUSH = io_store_cmd_payload_flush;
  assign store_pipeline_stages_0_FLUSH_FREE = io_store_cmd_payload_flushFree;
  assign store_pipeline_stages_0_PREFETCH = io_store_cmd_payload_prefetch;
  assign store_pipeline_stages_0_GENERATION = io_store_cmd_payload_generation;
  assign store_pipeline_stages_0_WAYS_HAZARD = 1'b0;
  assign io_store_cmd_ready = 1'b1;
  assign ways_0_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign ways_0_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[7 : 6];
  assign store_pipeline_stages_1_WAYS_TAGS_0_loaded = ways_0_storeRead_rsp_loaded;
  assign store_pipeline_stages_1_WAYS_TAGS_0_address = ways_0_storeRead_rsp_address;
  assign store_pipeline_stages_1_WAYS_TAGS_0_fault = ways_0_storeRead_rsp_fault;
  assign store_pipeline_stages_1_WAYS_HITS[0] = (store_pipeline_stages_1_WAYS_TAGS_0_loaded && (store_pipeline_stages_1_WAYS_TAGS_0_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 8]));
  assign store_pipeline_stages_1_WAYS_HIT = (|store_pipeline_stages_1_WAYS_HITS);
  assign status_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign status_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[7 : 6];
  assign store_pipeline_stages_1_STATUS_0_dirty = status_storeRead_rsp_0_dirty;
  always @(*) begin
    _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = store_pipeline_stages_1_STATUS_0_dirty;
    if(when_DataCache_l860_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = status_writeLast_payload_data_0_dirty;
    end
    if(when_DataCache_l863_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = status_write_payload_data_0_dirty;
    end
  end

  assign when_DataCache_l860_1 = (status_writeLast_valid && (status_writeLast_payload_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[7 : 6]));
  assign when_DataCache_l863_1 = (status_write_valid && (status_write_payload_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[7 : 6]));
  assign store_pipeline_stages_1_STATUS_overloaded_0_dirty = _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  always @(*) begin
    store_pipeline_stages_1_REFILL_HITS_EARLY = {(refill_slots_1_valid && (refill_slots_1_address[31 : 6] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 6])),(refill_slots_0_valid && (refill_slots_0_address[31 : 6] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 6]))};
    if(store_refillCheckEarly_refillPushHit) begin
      if(_zz_11) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[0] = 1'b1;
      end
      if(_zz_12) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[1] = 1'b1;
      end
    end
  end

  assign store_refillCheckEarly_refillPushHit = (refill_push_valid && (refill_push_payload_address[31 : 6] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 6]));
  assign store_pipeline_stages_2_REFILL_HITS = (store_pipeline_stages_2_REFILL_HITS_EARLY & {refill_slots_1_valid,refill_slots_0_valid});
  assign store_pipeline_stages_2_PROBE = 1'b0;
  always @(*) begin
    plru_fromStore_valid = 1'b0;
    if(store_ctrl_startRefill) begin
      plru_fromStore_valid = 1'b1;
    end
    if(store_ctrl_writeCache) begin
      plru_fromStore_valid = 1'b1;
    end
  end

  assign plru_fromStore_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 6];
  assign store_pipeline_stages_2_GENERATION_OK = (((store_pipeline_stages_2_GENERATION == store_target) || store_pipeline_stages_2_PREFETCH) || store_pipeline_stages_2_PROBE);
  always @(*) begin
    store_ctrl_reservation_take = 1'b0;
    if(when_DataCache_l1726) begin
      store_ctrl_reservation_take = 1'b1;
    end
  end

  assign store_ctrl_replacedWayNeedWriteback = (store_pipeline_stages_2_WAYS_TAGS_0_loaded && store_pipeline_stages_2_STATUS_0_dirty);
  assign store_ctrl_refillHit = (|(store_pipeline_stages_2_REFILL_HITS & {refill_slots_1_valid,refill_slots_0_valid}));
  assign store_ctrl_lineBusy = ((|{(refill_slots_1_valid && (refill_slots_1_address[7 : 6] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 6])),(refill_slots_0_valid && (refill_slots_0_address[7 : 6] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[7 : 6]))}) || 1'b0);
  assign store_ctrl_waysHitHazard = (|(store_pipeline_stages_2_WAYS_HITS & store_pipeline_stages_2_WAYS_HAZARD_resulting));
  assign store_ctrl_wasClean = (! (|(store_pipeline_stages_2_STATUS_0_dirty & store_pipeline_stages_2_WAYS_HITS)));
  assign store_ctrl_bankBusy = ((((! store_pipeline_stages_2_FLUSH) && (! store_pipeline_stages_2_PREFETCH)) && (! store_pipeline_stages_2_PROBE)) && (|(store_pipeline_stages_2_WAYS_HITS & refill_read_bankWriteNotif)));
  assign store_ctrl_hitUnique = 1'b1;
  assign store_ctrl_hitFault = (|(store_pipeline_stages_2_WAYS_HITS & store_pipeline_stages_2_WAYS_TAGS_0_fault));
  always @(*) begin
    store_pipeline_stages_2_REDO = (((((store_pipeline_stages_2_MISS || store_ctrl_waysHitHazard) || store_ctrl_bankBusy) || store_ctrl_refillHit) || (store_ctrl_wasClean && (! store_ctrl_reservation_win))) || (! store_ctrl_hitUnique));
    if(store_pipeline_stages_2_FLUSH) begin
      store_pipeline_stages_2_REDO = (store_ctrl_needFlush || (|store_pipeline_stages_2_WAYS_HAZARD_resulting));
    end
    if(store_pipeline_stages_2_IO) begin
      store_pipeline_stages_2_REDO = 1'b0;
    end
  end

  always @(*) begin
    store_pipeline_stages_2_MISS = (((! store_pipeline_stages_2_WAYS_HIT) && (! store_ctrl_waysHitHazard)) && (! store_ctrl_refillHit));
    if(store_pipeline_stages_2_IO) begin
      store_pipeline_stages_2_MISS = 1'b0;
    end
  end

  assign store_ctrl_canRefill = (((((! refill_full) && (! store_ctrl_lineBusy)) && (! load_ctrl_startRefill)) && store_ctrl_reservation_win) && (! store_pipeline_stages_2_WAYS_HAZARD_resulting[0]));
  assign store_ctrl_askRefill = (((store_pipeline_stages_2_MISS && store_ctrl_canRefill) && (! store_ctrl_refillHit)) && (! (store_ctrl_replacedWayNeedWriteback && writeback_full)));
  assign store_ctrl_askUpgrade = (((! store_pipeline_stages_2_MISS) && store_ctrl_canRefill) && (! store_ctrl_hitUnique));
  always @(*) begin
    store_ctrl_startRefill = ((store_pipeline_stages_2_valid && store_pipeline_stages_2_GENERATION_OK) && store_ctrl_askRefill);
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_startRefill = 1'b0;
    end
  end

  always @(*) begin
    store_ctrl_startUpgrade = ((store_pipeline_stages_2_valid && store_pipeline_stages_2_GENERATION_OK) && store_ctrl_askUpgrade);
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_startUpgrade = 1'b0;
    end
    if(store_pipeline_stages_2_IO) begin
      store_ctrl_startUpgrade = 1'b0;
    end
  end

  assign store_pipeline_stages_2_REFILL_SLOT_FULL = ((store_pipeline_stages_2_MISS && (! store_ctrl_refillHit)) && refill_full);
  assign store_pipeline_stages_2_REFILL_SLOT = ((store_ctrl_askRefill || store_ctrl_askUpgrade) ? refill_free : 2'b00);
  always @(*) begin
    store_ctrl_writeCache = ((((store_pipeline_stages_2_valid && store_pipeline_stages_2_GENERATION_OK) && (! store_pipeline_stages_2_REDO)) && (! store_pipeline_stages_2_PREFETCH)) && (! store_pipeline_stages_2_PROBE));
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_writeCache = 1'b0;
    end
    if(store_pipeline_stages_2_IO) begin
      store_ctrl_writeCache = 1'b0;
    end
  end

  always @(*) begin
    store_ctrl_setDirty = (store_ctrl_writeCache && store_ctrl_wasClean);
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_setDirty = 1'b0;
    end
    if(store_pipeline_stages_2_IO) begin
      store_ctrl_setDirty = 1'b0;
    end
  end

  assign store_ctrl_needFlushs = (store_pipeline_stages_2_WAYS_TAGS_0_loaded & store_pipeline_stages_2_STATUS_0_dirty);
  assign store_ctrl_needFlushs_bools_0 = store_ctrl_needFlushs[0];
  assign _zz_store_ctrl_needFlushOh[0] = (store_ctrl_needFlushs_bools_0 && (! 1'b0));
  assign store_ctrl_needFlushOh = _zz_store_ctrl_needFlushOh;
  assign _zz_15 = store_ctrl_needFlushOh[0];
  assign store_ctrl_needFlush = (|store_ctrl_needFlushs);
  assign store_ctrl_canFlush = (((store_ctrl_reservation_win && (! writeback_full)) && (! (|{refill_slots_1_valid,refill_slots_0_valid}))) && (! (|store_pipeline_stages_2_WAYS_HAZARD_resulting)));
  assign store_ctrl_startFlush = ((((store_pipeline_stages_2_valid && store_pipeline_stages_2_FLUSH) && store_pipeline_stages_2_GENERATION_OK) && store_ctrl_needFlush) && store_ctrl_canFlush);
  assign when_DataCache_l1726 = (((store_ctrl_startRefill || store_ctrl_startUpgrade) || store_ctrl_setDirty) || store_ctrl_startFlush);
  assign when_DataCache_l1733 = (store_ctrl_startRefill || store_ctrl_startFlush);
  assign when_DataCache_l1751 = (store_ctrl_startRefill || store_ctrl_startUpgrade);
  assign when_DataCache_l1775 = store_pipeline_stages_2_WAYS_HITS[0];
  assign when_DataCache_l1805 = ((((store_pipeline_stages_2_valid && store_pipeline_stages_2_REDO) && store_pipeline_stages_2_GENERATION_OK) && (! store_pipeline_stages_2_PREFETCH)) && (! store_pipeline_stages_2_PROBE));
  assign io_store_rsp_valid = (store_pipeline_stages_2_valid && (! store_pipeline_stages_2_PROBE));
  assign io_store_rsp_payload_generationKo = (! store_pipeline_stages_2_GENERATION_OK);
  assign io_store_rsp_payload_fault = 1'b0;
  assign io_store_rsp_payload_redo = store_pipeline_stages_2_REDO;
  assign io_store_rsp_payload_refillSlotAny = store_pipeline_stages_2_REFILL_SLOT_FULL;
  assign io_store_rsp_payload_refillSlot = store_pipeline_stages_2_REFILL_SLOT;
  assign io_store_rsp_payload_flush = store_pipeline_stages_2_FLUSH;
  assign io_store_rsp_payload_prefetch = store_pipeline_stages_2_PREFETCH;
  assign io_store_rsp_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  assign io_store_rsp_payload_io = store_pipeline_stages_2_IO;
  assign store_pipeline_stages_2_isThrown = store_pipeline_stages_2_throwRequest_DataCache_l1552;
  assign store_pipeline_stages_1_isThrown = store_pipeline_stages_1_throwRequest_DataCache_l1552;
  assign store_pipeline_stages_0_isThrown = store_pipeline_stages_0_throwRequest_DataCache_l1552;
  always @(*) begin
    _zz_store_pipeline_stages_1_valid = store_pipeline_stages_0_valid;
    if(when_Pipeline_l272_2) begin
      _zz_store_pipeline_stages_1_valid = 1'b0;
    end
  end

  assign when_Pipeline_l272_2 = (|store_pipeline_discardAll);
  always @(*) begin
    _zz_store_pipeline_stages_2_valid = store_pipeline_stages_1_valid;
    if(when_Pipeline_l272_3) begin
      _zz_store_pipeline_stages_2_valid = 1'b0;
    end
  end

  assign store_pipeline_stages_1_ready = 1'b1;
  assign when_Pipeline_l272_3 = (|store_pipeline_discardAll);
  assign store_pipeline_stages_2_WAYS_HAZARD_resulting = store_pipeline_stages_2_WAYS_HAZARD_overloaded;
  assign io_refillEvent = refill_push_valid;
  assign io_writebackEvent = writeback_push_valid;
  assign io_tagEvent = (|waysWrite_mask);
  assign invalidate_reservation_win = (! 1'b0);
  assign refill_read_reservation_win = (! 1'b0);
  assign load_ctrl_reservation_win = (! (|{refill_read_reservation_take,invalidate_reservation_take}));
  assign store_ctrl_reservation_win = (! (|{load_ctrl_reservation_take,{refill_read_reservation_take,invalidate_reservation_take}}));
  always @(posedge clk) begin
    waysWrite_maskLast <= waysWrite_mask;
    waysWrite_addressLast <= waysWrite_address;
    status_writeLast_payload_address <= status_write_payload_address;
    status_writeLast_payload_data_0_dirty <= status_write_payload_data_0_dirty;
    refill_slots_0_loadedCounter <= (refill_slots_0_loadedCounter + (refill_slots_0_loaded && (! refill_slots_0_loadedDone)));
    refill_slots_1_loadedCounter <= (refill_slots_1_loadedCounter + (refill_slots_1_loaded && (! refill_slots_1_loadedDone)));
    if(refill_push_valid) begin
      if(when_DataCache_l961) begin
        refill_slots_0_address <= refill_push_payload_address;
        refill_slots_0_cmdSent <= 1'b0;
        refill_slots_0_priority <= 1'b1;
        refill_slots_0_loaded <= 1'b0;
        refill_slots_0_loadedCounter <= 1'b0;
        refill_slots_0_victim <= refill_push_payload_victim;
        refill_slots_0_writebackHazards <= 2'b00;
      end else begin
        if(_zz_12) begin
          refill_slots_0_priority[0] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_DataCache_l961_1) begin
        refill_slots_1_address <= refill_push_payload_address;
        refill_slots_1_cmdSent <= 1'b0;
        refill_slots_1_priority <= 1'b1;
        refill_slots_1_loaded <= 1'b0;
        refill_slots_1_loadedCounter <= 1'b0;
        refill_slots_1_victim <= refill_push_payload_victim;
        refill_slots_1_writebackHazards <= 2'b00;
      end else begin
        if(_zz_11) begin
          refill_slots_1_priority[0] <= 1'b0;
        end
      end
    end
    if(refill_read_arbiter_oh[0]) begin
      refill_slots_0_writebackHazards <= refill_read_writebackHazards;
      if(when_DataCache_l998) begin
        refill_slots_0_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel) begin
      refill_slots_1_writebackHazards <= refill_read_writebackHazards;
      if(when_DataCache_l998_1) begin
        refill_slots_1_cmdSent <= 1'b1;
      end
    end
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1037) begin
        case(io_mem_read_rsp_payload_id)
          1'b0 : begin
            refill_slots_0_loaded <= 1'b1;
          end
          default : begin
            refill_slots_1_loaded <= 1'b1;
          end
        endcase
      end
    end
    if(writeback_slots_0_fire) begin
      refill_slots_0_writebackHazards[0] <= 1'b0;
      refill_slots_1_writebackHazards[0] <= 1'b0;
    end
    if(writeback_slots_1_fire) begin
      refill_slots_0_writebackHazards[1] <= 1'b0;
      refill_slots_1_writebackHazards[1] <= 1'b0;
    end
    if(writeback_push_valid) begin
      if(when_DataCache_l1128) begin
        writeback_slots_0_address <= writeback_push_payload_address;
        writeback_slots_0_writeCmdDone <= 1'b0;
        writeback_slots_0_priority <= 1'b1;
        writeback_slots_0_readCmdDone <= 1'b0;
        writeback_slots_0_readRspDone <= 1'b0;
        writeback_slots_0_victimBufferReady <= 1'b0;
      end else begin
        if(writeback_free[1]) begin
          writeback_slots_0_priority[0] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_DataCache_l1128_1) begin
        writeback_slots_1_address <= writeback_push_payload_address;
        writeback_slots_1_writeCmdDone <= 1'b0;
        writeback_slots_1_priority <= 1'b1;
        writeback_slots_1_readCmdDone <= 1'b0;
        writeback_slots_1_readRspDone <= 1'b0;
        writeback_slots_1_victimBufferReady <= 1'b0;
      end else begin
        if(writeback_free[0]) begin
          writeback_slots_1_priority[0] <= 1'b0;
        end
      end
    end
    if(when_DataCache_l1175) begin
      if(writeback_read_arbiter_oh[0]) begin
        writeback_slots_0_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel) begin
        writeback_slots_1_readCmdDone <= 1'b1;
      end
    end
    if(writeback_read_slotRead_valid) begin
      refill_slots_0_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_1_victim[writeback_read_slotRead_payload_id] <= 1'b0;
    end
    writeback_read_slotReadLast_payload_id <= writeback_read_slotRead_payload_id;
    writeback_read_slotReadLast_payload_last <= writeback_read_slotRead_payload_last;
    writeback_read_slotReadLast_payload_wordIndex <= writeback_read_slotRead_payload_wordIndex;
    if(writeback_read_slotReadLast_valid) begin
      case(writeback_read_slotReadLast_payload_id)
        1'b0 : begin
          writeback_slots_0_victimBufferReady <= 1'b1;
        end
        default : begin
          writeback_slots_1_victimBufferReady <= 1'b1;
        end
      endcase
      if(writeback_read_slotReadLast_payload_last) begin
        case(writeback_read_slotReadLast_payload_id)
          1'b0 : begin
            writeback_slots_0_readRspDone <= 1'b1;
          end
          default : begin
            writeback_slots_1_readRspDone <= 1'b1;
          end
        endcase
      end
    end
    if(when_DataCache_l1253) begin
      if(writeback_write_arbiter_oh[0]) begin
        writeback_slots_0_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel) begin
        writeback_slots_1_writeCmdDone <= 1'b1;
      end
    end
    if(writeback_write_bufferRead_ready) begin
      writeback_write_bufferRead_rData_id <= writeback_write_bufferRead_payload_id;
      writeback_write_bufferRead_rData_address <= writeback_write_bufferRead_payload_address;
      writeback_write_bufferRead_rData_last <= writeback_write_bufferRead_payload_last;
    end
    load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION <= load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION;
    load_pipeline_stages_1_WAYS_HAZARD <= load_pipeline_stages_0_WAYS_HAZARD;
    load_pipeline_stages_1_UNLOCKED <= load_pipeline_stages_0_UNLOCKED;
    load_pipeline_stages_1_NEED_UNIQUE <= load_pipeline_stages_0_NEED_UNIQUE;
    load_pipeline_stages_1_BANK_BUSY <= load_pipeline_stages_0_BANK_BUSY_overloaded;
    load_pipeline_stages_2_WAYS_HAZARD <= load_pipeline_stages_1_WAYS_HAZARD_overloaded;
    load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION <= load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION;
    load_pipeline_stages_2_BANK_BUSY_REMAPPED <= load_pipeline_stages_1_BANK_BUSY_REMAPPED;
    load_pipeline_stages_2_BANKS_MUXES_0 <= load_pipeline_stages_1_BANKS_MUXES_0;
    load_pipeline_stages_2_ADDRESS_POST_TRANSLATION <= load_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
    load_pipeline_stages_2_ABORD <= load_pipeline_stages_1_ABORD;
    load_pipeline_stages_2_WAYS_TAGS_0_loaded <= load_pipeline_stages_1_WAYS_TAGS_0_loaded;
    load_pipeline_stages_2_WAYS_TAGS_0_address <= load_pipeline_stages_1_WAYS_TAGS_0_address;
    load_pipeline_stages_2_WAYS_TAGS_0_fault <= load_pipeline_stages_1_WAYS_TAGS_0_fault;
    load_pipeline_stages_2_WAYS_HITS <= load_pipeline_stages_1_WAYS_HITS;
    load_pipeline_stages_2_STATUS_0_dirty <= load_pipeline_stages_1_STATUS_overloaded_0_dirty;
    load_pipeline_stages_2_LOCKED <= load_pipeline_stages_1_LOCKED;
    load_pipeline_stages_2_NEED_UNIQUE <= load_pipeline_stages_1_NEED_UNIQUE;
    store_pipeline_stages_1_ADDRESS_POST_TRANSLATION <= store_pipeline_stages_0_ADDRESS_POST_TRANSLATION;
    store_pipeline_stages_1_CPU_WORD <= store_pipeline_stages_0_CPU_WORD;
    store_pipeline_stages_1_CPU_MASK <= store_pipeline_stages_0_CPU_MASK;
    store_pipeline_stages_1_IO <= store_pipeline_stages_0_IO;
    store_pipeline_stages_1_FLUSH <= store_pipeline_stages_0_FLUSH;
    store_pipeline_stages_1_FLUSH_FREE <= store_pipeline_stages_0_FLUSH_FREE;
    store_pipeline_stages_1_PREFETCH <= store_pipeline_stages_0_PREFETCH;
    store_pipeline_stages_1_GENERATION <= store_pipeline_stages_0_GENERATION;
    store_pipeline_stages_1_WAYS_HAZARD <= store_pipeline_stages_0_WAYS_HAZARD;
    store_pipeline_stages_2_WAYS_HAZARD <= store_pipeline_stages_1_WAYS_HAZARD_overloaded;
    store_pipeline_stages_2_ADDRESS_POST_TRANSLATION <= store_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
    store_pipeline_stages_2_WAYS_TAGS_0_loaded <= store_pipeline_stages_1_WAYS_TAGS_0_loaded;
    store_pipeline_stages_2_WAYS_TAGS_0_address <= store_pipeline_stages_1_WAYS_TAGS_0_address;
    store_pipeline_stages_2_WAYS_TAGS_0_fault <= store_pipeline_stages_1_WAYS_TAGS_0_fault;
    store_pipeline_stages_2_WAYS_HITS <= store_pipeline_stages_1_WAYS_HITS;
    store_pipeline_stages_2_WAYS_HIT <= store_pipeline_stages_1_WAYS_HIT;
    store_pipeline_stages_2_STATUS_0_dirty <= store_pipeline_stages_1_STATUS_overloaded_0_dirty;
    store_pipeline_stages_2_REFILL_HITS_EARLY <= store_pipeline_stages_1_REFILL_HITS_EARLY;
    store_pipeline_stages_2_GENERATION <= store_pipeline_stages_1_GENERATION;
    store_pipeline_stages_2_PREFETCH <= store_pipeline_stages_1_PREFETCH;
    store_pipeline_stages_2_FLUSH <= store_pipeline_stages_1_FLUSH;
    store_pipeline_stages_2_IO <= store_pipeline_stages_1_IO;
    store_pipeline_stages_2_CPU_WORD <= store_pipeline_stages_1_CPU_WORD;
    store_pipeline_stages_2_CPU_MASK <= store_pipeline_stages_1_CPU_MASK;
    store_pipeline_stages_2_FLUSH_FREE <= store_pipeline_stages_1_FLUSH_FREE;
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      status_writeLast_valid <= 1'b0;
      invalidate_counter <= 3'b000;
      invalidate_firstEver <= 1'b1;
      refill_slots_0_valid <= 1'b0;
      refill_slots_1_valid <= 1'b0;
      refill_pushCounter <= 32'h00000000;
      refill_read_arbiter_lock <= 2'b00;
      refill_read_wordIndex <= 4'b0000;
      refill_read_hadError <= 1'b0;
      writeback_slots_0_valid <= 1'b0;
      writeback_slots_1_valid <= 1'b0;
      writeback_read_arbiter_lock <= 2'b00;
      writeback_read_wordIndex <= 4'b0000;
      writeback_read_slotReadLast_valid <= 1'b0;
      writeback_write_arbiter_lock <= 2'b00;
      writeback_write_wordIndex <= 4'b0000;
      writeback_write_bufferRead_rValid <= 1'b0;
      load_pipeline_stages_1_valid <= 1'b0;
      load_pipeline_stages_2_valid <= 1'b0;
      store_target <= 1'b0;
      store_pipeline_stages_1_valid <= 1'b0;
      store_pipeline_stages_2_valid <= 1'b0;
    end else begin
      status_writeLast_valid <= status_write_valid;
      if(when_DataCache_l888) begin
        invalidate_counter <= (invalidate_counter + 3'b001);
      end
      if(invalidate_done) begin
        invalidate_firstEver <= 1'b0;
      end
      if(when_DataCache_l934) begin
        refill_slots_0_valid <= 1'b0;
      end
      if(when_DataCache_l934_1) begin
        refill_slots_1_valid <= 1'b0;
      end
      if(refill_push_valid) begin
        refill_pushCounter <= (refill_pushCounter + 32'h00000001);
      end
      if(refill_push_valid) begin
        if(when_DataCache_l961) begin
          refill_slots_0_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_DataCache_l961_1) begin
          refill_slots_1_valid <= 1'b1;
        end
      end
      refill_read_arbiter_lock <= refill_read_arbiter_oh;
      if(when_DataCache_l986) begin
        refill_read_arbiter_lock <= 2'b00;
      end
      if(when_DataCache_l1026) begin
        refill_read_hadError <= 1'b1;
      end
      if(io_mem_read_rsp_valid) begin
        if(refill_read_rspWithData) begin
          refill_read_wordIndex <= (refill_read_wordIndex + 4'b0001);
        end
        if(when_DataCache_l1037) begin
          refill_read_hadError <= 1'b0;
        end
      end
      if(writeback_slots_0_fire) begin
        writeback_slots_0_valid <= 1'b0;
      end
      if(writeback_slots_1_fire) begin
        writeback_slots_1_valid <= 1'b0;
      end
      if(writeback_push_valid) begin
        if(when_DataCache_l1128) begin
          writeback_slots_0_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_DataCache_l1128_1) begin
          writeback_slots_1_valid <= 1'b1;
        end
      end
      writeback_read_arbiter_lock <= writeback_read_arbiter_oh;
      writeback_read_wordIndex <= (writeback_read_wordIndex + _zz_writeback_read_wordIndex);
      if(when_DataCache_l1175) begin
        writeback_read_arbiter_lock <= 2'b00;
      end
      writeback_read_slotReadLast_valid <= writeback_read_slotRead_valid;
      writeback_write_arbiter_lock <= writeback_write_arbiter_oh;
      writeback_write_wordIndex <= (writeback_write_wordIndex + _zz_writeback_write_wordIndex);
      if(when_DataCache_l1253) begin
        writeback_write_arbiter_lock <= 2'b00;
      end
      if(writeback_write_bufferRead_ready) begin
        writeback_write_bufferRead_rValid <= writeback_write_bufferRead_valid;
      end
      load_pipeline_stages_1_valid <= _zz_load_pipeline_stages_1_valid;
      load_pipeline_stages_2_valid <= _zz_load_pipeline_stages_2_valid;
      if(when_DataCache_l1805) begin
        store_target <= (! store_target);
      end
      store_pipeline_stages_1_valid <= _zz_store_pipeline_stages_1_valid;
      store_pipeline_stages_2_valid <= _zz_store_pipeline_stages_2_valid;
    end
  end


endmodule

module AllocatorMultiPortMem (
  input  wire          io_push_0_valid /* verilator public */ ,
  input  wire [5:0]    io_push_0_payload /* verilator public */ ,
  input  wire [0:0]    io_pop_mask /* verilator public */ ,
  output wire          io_pop_ready /* verilator public */ ,
  input  wire          io_pop_fire /* verilator public */ ,
  output wire [5:0]    io_pop_values_0 /* verilator public */ ,
  input  wire          clk,
  input  wire          reset
);

  wire       [5:0]    ways_0_mem_spinal_port1;
  reg        [0:0]    _zz_popMaskCount;
  wire       [0:0]    _zz_popMaskCount_1;
  reg        [0:0]    _zz_ptr_pushCount;
  wire       [0:0]    _zz_ptr_pushCount_1;
  wire       [6:0]    _zz_ptr_push;
  wire       [6:0]    _zz_ptr_pop;
  wire       [6:0]    _zz_ptr_occupancy;
  wire       [6:0]    _zz_ptr_occupancy_1;
  wire       [6:0]    _zz_ptr_occupancy_2;
  wire       [0:0]    _zz_ptr_occupancy_3;
  wire       [6:0]    _zz_pushArbitration_pushOffset_1;
  wire       [0:0]    _zz_pushArbitration_pushOffset_1_1;
  wire       [5:0]    _zz_ways_0_mem_port;
  wire       [5:0]    _zz_ways_0_mem_port_1;
  wire                _zz_ways_0_mem_port_2;
  wire       [6:0]    _zz_popArbitration_popOffset_1;
  wire       [0:0]    _zz_popArbitration_popOffset_1_1;
  reg        [6:0]    popArbitration_popOffset_1;
  reg        [6:0]    pushArbitration_pushOffset_1;
  wire       [0:0]    popMaskCount;
  reg        [6:0]    ptr_push;
  reg        [6:0]    ptr_pop;
  reg        [6:0]    ptr_occupancy;
  wire       [0:0]    ptr_pushCount;
  wire       [6:0]    pushArbitration_pushOffset;
  wire       [6:0]    pushArbitration_push_0_ptr;
  wire       [6:0]    ways_0_push_offset;
  wire       [0:0]    ways_0_push_hits;
  wire       [6:0]    ways_0_pop_offset;
  wire       [5:0]    _zz_ways_0_pop_data;
  wire       [5:0]    ways_0_pop_data;
  wire       [6:0]    popArbitration_popOffset;
  wire       [6:0]    popArbitration_pop_0_ptr;
  (* ram_style = "distributed" *) reg [5:0] ways_0_mem [0:63];

  assign _zz_ptr_push = {6'd0, ptr_pushCount};
  assign _zz_ptr_pop = {6'd0, popMaskCount};
  assign _zz_ptr_occupancy = (ptr_occupancy + _zz_ptr_occupancy_1);
  assign _zz_ptr_occupancy_1 = {6'd0, ptr_pushCount};
  assign _zz_ptr_occupancy_3 = (io_pop_fire ? popMaskCount : 1'b0);
  assign _zz_ptr_occupancy_2 = {6'd0, _zz_ptr_occupancy_3};
  assign _zz_pushArbitration_pushOffset_1_1 = io_push_0_valid;
  assign _zz_pushArbitration_pushOffset_1 = {6'd0, _zz_pushArbitration_pushOffset_1_1};
  assign _zz_popArbitration_popOffset_1_1 = io_pop_mask[0];
  assign _zz_popArbitration_popOffset_1 = {6'd0, _zz_popArbitration_popOffset_1_1};
  assign _zz_ways_0_mem_port = ways_0_push_offset[5 : 0];
  assign _zz_ways_0_mem_port_1 = io_push_0_payload;
  assign _zz_ways_0_mem_port_2 = (|ways_0_push_hits);
  assign _zz_popMaskCount_1 = io_pop_mask[0];
  assign _zz_ptr_pushCount_1 = io_push_0_valid;
  always @(posedge clk) begin
    if(_zz_ways_0_mem_port_2) begin
      ways_0_mem[_zz_ways_0_mem_port] <= _zz_ways_0_mem_port_1;
    end
  end

  assign ways_0_mem_spinal_port1 = ways_0_mem[_zz_ways_0_pop_data];
  always @(*) begin
    case(_zz_popMaskCount_1)
      1'b0 : _zz_popMaskCount = 1'b0;
      default : _zz_popMaskCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_ptr_pushCount_1)
      1'b0 : _zz_ptr_pushCount = 1'b0;
      default : _zz_ptr_pushCount = 1'b1;
    endcase
  end

  always @(*) begin
    popArbitration_popOffset_1 = popArbitration_popOffset;
    popArbitration_popOffset_1 = (popArbitration_popOffset + _zz_popArbitration_popOffset_1);
  end

  always @(*) begin
    pushArbitration_pushOffset_1 = pushArbitration_pushOffset;
    pushArbitration_pushOffset_1 = (pushArbitration_pushOffset + _zz_pushArbitration_pushOffset_1);
  end

  assign popMaskCount = _zz_popMaskCount;
  assign ptr_pushCount = _zz_ptr_pushCount;
  assign pushArbitration_pushOffset = ptr_push;
  assign pushArbitration_push_0_ptr = pushArbitration_pushOffset;
  assign ways_0_push_offset = (ptr_push + 7'h00);
  assign ways_0_push_hits = (io_push_0_valid & 1'b1);
  assign ways_0_pop_offset = (ptr_pop + 7'h00);
  assign _zz_ways_0_pop_data = ways_0_pop_offset[5 : 0];
  assign ways_0_pop_data = ways_0_mem_spinal_port1;
  assign popArbitration_popOffset = ptr_pop;
  assign popArbitration_pop_0_ptr = popArbitration_popOffset;
  assign io_pop_values_0 = ways_0_pop_data;
  assign io_pop_ready = (7'h01 <= ptr_occupancy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      ptr_push <= 7'h00;
      ptr_pop <= 7'h00;
      ptr_occupancy <= 7'h00;
    end else begin
      ptr_push <= (ptr_push + _zz_ptr_push);
      if(io_pop_fire) begin
        ptr_pop <= (ptr_pop + _zz_ptr_pop);
      end
      ptr_occupancy <= (_zz_ptr_occupancy - _zz_ptr_occupancy_2);
    end
  end


endmodule

module TranslatorWithRollback (
  input  wire          io_rollback,
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_payload_address,
  input  wire [5:0]    io_writes_0_payload_data,
  input  wire          io_commits_0_valid,
  input  wire [4:0]    io_commits_0_payload_address,
  input  wire [5:0]    io_commits_0_payload_data,
  input  wire          io_reads_0_cmd_valid,
  input  wire [4:0]    io_reads_0_cmd_payload,
  output wire          io_reads_0_rsp_valid,
  output wire [5:0]    io_reads_0_rsp_payload,
  input  wire          io_reads_1_cmd_valid,
  input  wire [4:0]    io_reads_1_cmd_payload,
  output wire          io_reads_1_rsp_valid,
  output wire [5:0]    io_reads_1_rsp_payload,
  input  wire          io_reads_2_cmd_valid,
  input  wire [4:0]    io_reads_2_cmd_payload,
  output wire          io_reads_2_rsp_valid,
  output wire [5:0]    io_reads_2_rsp_payload,
  input  wire          clk,
  input  wire          reset
);

  wire       [5:0]    writes_ram_spinal_port1;
  wire       [5:0]    writes_ram_spinal_port2;
  wire       [5:0]    writes_ram_spinal_port3;
  wire       [5:0]    commits_ram_spinal_port1;
  wire       [5:0]    commits_ram_spinal_port2;
  wire       [5:0]    commits_ram_spinal_port3;
  wire       [5:0]    _zz_writes_ram_port;
  wire                _zz_writes_ram_port_1;
  wire       [5:0]    _zz_commits_ram_port;
  wire                _zz_commits_ram_port_1;
  reg        [31:0]   location_updated;
  wire                location_set_0_hits_0;
  wire                when_RfTranslationPlugin_l71;
  wire                location_set_1_hits_0;
  wire                when_RfTranslationPlugin_l71_1;
  wire                location_set_2_hits_0;
  wire                when_RfTranslationPlugin_l71_2;
  wire                location_set_3_hits_0;
  wire                when_RfTranslationPlugin_l71_3;
  wire                location_set_4_hits_0;
  wire                when_RfTranslationPlugin_l71_4;
  wire                location_set_5_hits_0;
  wire                when_RfTranslationPlugin_l71_5;
  wire                location_set_6_hits_0;
  wire                when_RfTranslationPlugin_l71_6;
  wire                location_set_7_hits_0;
  wire                when_RfTranslationPlugin_l71_7;
  wire                location_set_8_hits_0;
  wire                when_RfTranslationPlugin_l71_8;
  wire                location_set_9_hits_0;
  wire                when_RfTranslationPlugin_l71_9;
  wire                location_set_10_hits_0;
  wire                when_RfTranslationPlugin_l71_10;
  wire                location_set_11_hits_0;
  wire                when_RfTranslationPlugin_l71_11;
  wire                location_set_12_hits_0;
  wire                when_RfTranslationPlugin_l71_12;
  wire                location_set_13_hits_0;
  wire                when_RfTranslationPlugin_l71_13;
  wire                location_set_14_hits_0;
  wire                when_RfTranslationPlugin_l71_14;
  wire                location_set_15_hits_0;
  wire                when_RfTranslationPlugin_l71_15;
  wire                location_set_16_hits_0;
  wire                when_RfTranslationPlugin_l71_16;
  wire                location_set_17_hits_0;
  wire                when_RfTranslationPlugin_l71_17;
  wire                location_set_18_hits_0;
  wire                when_RfTranslationPlugin_l71_18;
  wire                location_set_19_hits_0;
  wire                when_RfTranslationPlugin_l71_19;
  wire                location_set_20_hits_0;
  wire                when_RfTranslationPlugin_l71_20;
  wire                location_set_21_hits_0;
  wire                when_RfTranslationPlugin_l71_21;
  wire                location_set_22_hits_0;
  wire                when_RfTranslationPlugin_l71_22;
  wire                location_set_23_hits_0;
  wire                when_RfTranslationPlugin_l71_23;
  wire                location_set_24_hits_0;
  wire                when_RfTranslationPlugin_l71_24;
  wire                location_set_25_hits_0;
  wire                when_RfTranslationPlugin_l71_25;
  wire                location_set_26_hits_0;
  wire                when_RfTranslationPlugin_l71_26;
  wire                location_set_27_hits_0;
  wire                when_RfTranslationPlugin_l71_27;
  wire                location_set_28_hits_0;
  wire                when_RfTranslationPlugin_l71_28;
  wire                location_set_29_hits_0;
  wire                when_RfTranslationPlugin_l71_29;
  wire                location_set_30_hits_0;
  wire                when_RfTranslationPlugin_l71_30;
  wire                location_set_31_hits_0;
  wire                when_RfTranslationPlugin_l71_31;
  wire       [5:0]    read_0_written;
  wire       [5:0]    read_0_commited;
  wire                read_0_sel;
  wire       [5:0]    read_0_muxed;
  wire       [5:0]    read_1_written;
  wire       [5:0]    read_1_commited;
  wire                read_1_sel;
  wire       [5:0]    read_1_muxed;
  wire       [5:0]    read_2_written;
  wire       [5:0]    read_2_commited;
  wire                read_2_sel;
  wire       [5:0]    read_2_muxed;
  (* ram_style = "distributed" *) reg [5:0] writes_ram [0:31];
  (* ram_style = "distributed" *) reg [5:0] commits_ram [0:31];

  assign _zz_writes_ram_port = io_writes_0_payload_data;
  assign _zz_writes_ram_port_1 = (io_writes_0_valid && (! 1'b0));
  assign _zz_commits_ram_port = io_commits_0_payload_data;
  assign _zz_commits_ram_port_1 = (io_commits_0_valid && (! 1'b0));
  always @(posedge clk) begin
    if(_zz_writes_ram_port_1) begin
      writes_ram[io_writes_0_payload_address] <= _zz_writes_ram_port;
    end
  end

  assign writes_ram_spinal_port1 = writes_ram[io_reads_0_cmd_payload];
  assign writes_ram_spinal_port2 = writes_ram[io_reads_1_cmd_payload];
  assign writes_ram_spinal_port3 = writes_ram[io_reads_2_cmd_payload];
  always @(posedge clk) begin
    if(_zz_commits_ram_port_1) begin
      commits_ram[io_commits_0_payload_address] <= _zz_commits_ram_port;
    end
  end

  assign commits_ram_spinal_port1 = commits_ram[io_reads_0_cmd_payload];
  assign commits_ram_spinal_port2 = commits_ram[io_reads_1_cmd_payload];
  assign commits_ram_spinal_port3 = commits_ram[io_reads_2_cmd_payload];
  assign location_set_0_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h00));
  assign when_RfTranslationPlugin_l71 = (|location_set_0_hits_0);
  assign location_set_1_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h01));
  assign when_RfTranslationPlugin_l71_1 = (|location_set_1_hits_0);
  assign location_set_2_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h02));
  assign when_RfTranslationPlugin_l71_2 = (|location_set_2_hits_0);
  assign location_set_3_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h03));
  assign when_RfTranslationPlugin_l71_3 = (|location_set_3_hits_0);
  assign location_set_4_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h04));
  assign when_RfTranslationPlugin_l71_4 = (|location_set_4_hits_0);
  assign location_set_5_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h05));
  assign when_RfTranslationPlugin_l71_5 = (|location_set_5_hits_0);
  assign location_set_6_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h06));
  assign when_RfTranslationPlugin_l71_6 = (|location_set_6_hits_0);
  assign location_set_7_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h07));
  assign when_RfTranslationPlugin_l71_7 = (|location_set_7_hits_0);
  assign location_set_8_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h08));
  assign when_RfTranslationPlugin_l71_8 = (|location_set_8_hits_0);
  assign location_set_9_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h09));
  assign when_RfTranslationPlugin_l71_9 = (|location_set_9_hits_0);
  assign location_set_10_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0a));
  assign when_RfTranslationPlugin_l71_10 = (|location_set_10_hits_0);
  assign location_set_11_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0b));
  assign when_RfTranslationPlugin_l71_11 = (|location_set_11_hits_0);
  assign location_set_12_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0c));
  assign when_RfTranslationPlugin_l71_12 = (|location_set_12_hits_0);
  assign location_set_13_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0d));
  assign when_RfTranslationPlugin_l71_13 = (|location_set_13_hits_0);
  assign location_set_14_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0e));
  assign when_RfTranslationPlugin_l71_14 = (|location_set_14_hits_0);
  assign location_set_15_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0f));
  assign when_RfTranslationPlugin_l71_15 = (|location_set_15_hits_0);
  assign location_set_16_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h10));
  assign when_RfTranslationPlugin_l71_16 = (|location_set_16_hits_0);
  assign location_set_17_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h11));
  assign when_RfTranslationPlugin_l71_17 = (|location_set_17_hits_0);
  assign location_set_18_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h12));
  assign when_RfTranslationPlugin_l71_18 = (|location_set_18_hits_0);
  assign location_set_19_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h13));
  assign when_RfTranslationPlugin_l71_19 = (|location_set_19_hits_0);
  assign location_set_20_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h14));
  assign when_RfTranslationPlugin_l71_20 = (|location_set_20_hits_0);
  assign location_set_21_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h15));
  assign when_RfTranslationPlugin_l71_21 = (|location_set_21_hits_0);
  assign location_set_22_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h16));
  assign when_RfTranslationPlugin_l71_22 = (|location_set_22_hits_0);
  assign location_set_23_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h17));
  assign when_RfTranslationPlugin_l71_23 = (|location_set_23_hits_0);
  assign location_set_24_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h18));
  assign when_RfTranslationPlugin_l71_24 = (|location_set_24_hits_0);
  assign location_set_25_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h19));
  assign when_RfTranslationPlugin_l71_25 = (|location_set_25_hits_0);
  assign location_set_26_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1a));
  assign when_RfTranslationPlugin_l71_26 = (|location_set_26_hits_0);
  assign location_set_27_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1b));
  assign when_RfTranslationPlugin_l71_27 = (|location_set_27_hits_0);
  assign location_set_28_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1c));
  assign when_RfTranslationPlugin_l71_28 = (|location_set_28_hits_0);
  assign location_set_29_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1d));
  assign when_RfTranslationPlugin_l71_29 = (|location_set_29_hits_0);
  assign location_set_30_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1e));
  assign when_RfTranslationPlugin_l71_30 = (|location_set_30_hits_0);
  assign location_set_31_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1f));
  assign when_RfTranslationPlugin_l71_31 = (|location_set_31_hits_0);
  assign read_0_written = writes_ram_spinal_port1;
  assign read_0_commited = commits_ram_spinal_port1;
  assign read_0_sel = location_updated[io_reads_0_cmd_payload];
  assign read_0_muxed = (read_0_sel ? read_0_written : read_0_commited);
  assign io_reads_0_rsp_valid = io_reads_0_cmd_valid;
  assign io_reads_0_rsp_payload = read_0_muxed;
  assign read_1_written = writes_ram_spinal_port2;
  assign read_1_commited = commits_ram_spinal_port2;
  assign read_1_sel = location_updated[io_reads_1_cmd_payload];
  assign read_1_muxed = (read_1_sel ? read_1_written : read_1_commited);
  assign io_reads_1_rsp_valid = io_reads_1_cmd_valid;
  assign io_reads_1_rsp_payload = read_1_muxed;
  assign read_2_written = writes_ram_spinal_port3;
  assign read_2_commited = commits_ram_spinal_port3;
  assign read_2_sel = location_updated[io_reads_2_cmd_payload];
  assign read_2_muxed = (read_2_sel ? read_2_written : read_2_commited);
  assign io_reads_2_rsp_valid = io_reads_2_cmd_valid;
  assign io_reads_2_rsp_payload = read_2_muxed;
  always @(posedge clk) begin
    if(when_RfTranslationPlugin_l71) begin
      location_updated[0] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_1) begin
      location_updated[1] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_2) begin
      location_updated[2] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_3) begin
      location_updated[3] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_4) begin
      location_updated[4] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_5) begin
      location_updated[5] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_6) begin
      location_updated[6] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_7) begin
      location_updated[7] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_8) begin
      location_updated[8] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_9) begin
      location_updated[9] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_10) begin
      location_updated[10] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_11) begin
      location_updated[11] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_12) begin
      location_updated[12] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_13) begin
      location_updated[13] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_14) begin
      location_updated[14] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_15) begin
      location_updated[15] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_16) begin
      location_updated[16] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_17) begin
      location_updated[17] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_18) begin
      location_updated[18] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_19) begin
      location_updated[19] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_20) begin
      location_updated[20] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_21) begin
      location_updated[21] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_22) begin
      location_updated[22] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_23) begin
      location_updated[23] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_24) begin
      location_updated[24] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_25) begin
      location_updated[25] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_26) begin
      location_updated[26] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_27) begin
      location_updated[27] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_28) begin
      location_updated[28] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_29) begin
      location_updated[29] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_30) begin
      location_updated[30] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_31) begin
      location_updated[31] <= 1'b1;
    end
    if(io_rollback) begin
      location_updated <= 32'h00000000;
    end
  end


endmodule

module AxiLite4Plic (
  input  wire          io_bus_aw_valid,
  output wire          io_bus_aw_ready,
  input  wire [21:0]   io_bus_aw_payload_addr,
  input  wire [2:0]    io_bus_aw_payload_prot,
  input  wire          io_bus_w_valid,
  output wire          io_bus_w_ready,
  input  wire [31:0]   io_bus_w_payload_data,
  input  wire [3:0]    io_bus_w_payload_strb,
  output wire          io_bus_b_valid,
  input  wire          io_bus_b_ready,
  output wire [1:0]    io_bus_b_payload_resp,
  input  wire          io_bus_ar_valid,
  output wire          io_bus_ar_ready,
  input  wire [21:0]   io_bus_ar_payload_addr,
  input  wire [2:0]    io_bus_ar_payload_prot,
  output wire          io_bus_r_valid,
  input  wire          io_bus_r_ready,
  output wire [31:0]   io_bus_r_payload_data,
  output wire [1:0]    io_bus_r_payload_resp,
  input  wire [30:0]   io_sources,
  output wire [1:0]    io_targets,
  input  wire          clk,
  input  wire          reset
);

  wire       [4:0]    _zz_targets_0_bestRequest_id_82;
  wire       [4:0]    _zz_targets_0_bestRequest_id_83;
  wire       [4:0]    _zz_targets_0_bestRequest_id_84;
  wire       [4:0]    _zz_targets_0_bestRequest_id_85;
  wire       [4:0]    _zz_targets_0_bestRequest_id_86;
  wire       [4:0]    _zz_targets_0_bestRequest_id_87;
  wire       [4:0]    _zz_targets_0_bestRequest_id_88;
  wire       [4:0]    _zz_targets_0_bestRequest_id_89;
  wire       [4:0]    _zz_targets_0_bestRequest_id_90;
  wire       [4:0]    _zz_targets_0_bestRequest_id_91;
  wire       [4:0]    _zz_targets_0_bestRequest_id_92;
  wire       [4:0]    _zz_targets_0_bestRequest_id_93;
  wire       [4:0]    _zz_targets_0_bestRequest_id_94;
  wire       [4:0]    _zz_targets_0_bestRequest_id_95;
  wire       [4:0]    _zz_targets_0_bestRequest_id_96;
  wire       [4:0]    _zz_targets_0_bestRequest_id_97;
  wire       [4:0]    _zz_targets_1_bestRequest_id_82;
  wire       [4:0]    _zz_targets_1_bestRequest_id_83;
  wire       [4:0]    _zz_targets_1_bestRequest_id_84;
  wire       [4:0]    _zz_targets_1_bestRequest_id_85;
  wire       [4:0]    _zz_targets_1_bestRequest_id_86;
  wire       [4:0]    _zz_targets_1_bestRequest_id_87;
  wire       [4:0]    _zz_targets_1_bestRequest_id_88;
  wire       [4:0]    _zz_targets_1_bestRequest_id_89;
  wire       [4:0]    _zz_targets_1_bestRequest_id_90;
  wire       [4:0]    _zz_targets_1_bestRequest_id_91;
  wire       [4:0]    _zz_targets_1_bestRequest_id_92;
  wire       [4:0]    _zz_targets_1_bestRequest_id_93;
  wire       [4:0]    _zz_targets_1_bestRequest_id_94;
  wire       [4:0]    _zz_targets_1_bestRequest_id_95;
  wire       [4:0]    _zz_targets_1_bestRequest_id_96;
  wire       [4:0]    _zz_targets_1_bestRequest_id_97;
  wire                _zz_gateways_0_ip;
  wire                _zz_gateways_1_ip;
  wire                _zz_gateways_2_ip;
  wire                _zz_gateways_3_ip;
  wire                _zz_gateways_4_ip;
  wire                _zz_gateways_5_ip;
  wire                _zz_gateways_6_ip;
  wire                _zz_gateways_7_ip;
  wire                _zz_gateways_8_ip;
  wire                _zz_gateways_9_ip;
  wire                _zz_gateways_10_ip;
  wire                _zz_gateways_11_ip;
  wire                _zz_gateways_12_ip;
  wire                _zz_gateways_13_ip;
  wire                _zz_gateways_14_ip;
  wire                _zz_gateways_15_ip;
  wire                _zz_gateways_16_ip;
  wire                _zz_gateways_17_ip;
  wire                _zz_gateways_18_ip;
  wire                _zz_gateways_19_ip;
  wire                _zz_gateways_20_ip;
  wire                _zz_gateways_21_ip;
  wire                _zz_gateways_22_ip;
  wire                _zz_gateways_23_ip;
  wire                _zz_gateways_24_ip;
  wire                _zz_gateways_25_ip;
  wire                _zz_gateways_26_ip;
  wire                _zz_gateways_27_ip;
  wire                _zz_gateways_28_ip;
  wire                _zz_gateways_29_ip;
  wire                _zz_gateways_30_ip;
  wire       [1:0]    gateways_0_priority;
  reg                 gateways_0_ip;
  reg                 gateways_0_waitCompletion;
  wire                when_PlicGateway_l21;
  wire       [1:0]    gateways_1_priority;
  reg                 gateways_1_ip;
  reg                 gateways_1_waitCompletion;
  wire                when_PlicGateway_l21_1;
  wire       [1:0]    gateways_2_priority;
  reg                 gateways_2_ip;
  reg                 gateways_2_waitCompletion;
  wire                when_PlicGateway_l21_2;
  wire       [1:0]    gateways_3_priority;
  reg                 gateways_3_ip;
  reg                 gateways_3_waitCompletion;
  wire                when_PlicGateway_l21_3;
  wire       [1:0]    gateways_4_priority;
  reg                 gateways_4_ip;
  reg                 gateways_4_waitCompletion;
  wire                when_PlicGateway_l21_4;
  wire       [1:0]    gateways_5_priority;
  reg                 gateways_5_ip;
  reg                 gateways_5_waitCompletion;
  wire                when_PlicGateway_l21_5;
  wire       [1:0]    gateways_6_priority;
  reg                 gateways_6_ip;
  reg                 gateways_6_waitCompletion;
  wire                when_PlicGateway_l21_6;
  wire       [1:0]    gateways_7_priority;
  reg                 gateways_7_ip;
  reg                 gateways_7_waitCompletion;
  wire                when_PlicGateway_l21_7;
  wire       [1:0]    gateways_8_priority;
  reg                 gateways_8_ip;
  reg                 gateways_8_waitCompletion;
  wire                when_PlicGateway_l21_8;
  wire       [1:0]    gateways_9_priority;
  reg                 gateways_9_ip;
  reg                 gateways_9_waitCompletion;
  wire                when_PlicGateway_l21_9;
  wire       [1:0]    gateways_10_priority;
  reg                 gateways_10_ip;
  reg                 gateways_10_waitCompletion;
  wire                when_PlicGateway_l21_10;
  wire       [1:0]    gateways_11_priority;
  reg                 gateways_11_ip;
  reg                 gateways_11_waitCompletion;
  wire                when_PlicGateway_l21_11;
  wire       [1:0]    gateways_12_priority;
  reg                 gateways_12_ip;
  reg                 gateways_12_waitCompletion;
  wire                when_PlicGateway_l21_12;
  wire       [1:0]    gateways_13_priority;
  reg                 gateways_13_ip;
  reg                 gateways_13_waitCompletion;
  wire                when_PlicGateway_l21_13;
  wire       [1:0]    gateways_14_priority;
  reg                 gateways_14_ip;
  reg                 gateways_14_waitCompletion;
  wire                when_PlicGateway_l21_14;
  wire       [1:0]    gateways_15_priority;
  reg                 gateways_15_ip;
  reg                 gateways_15_waitCompletion;
  wire                when_PlicGateway_l21_15;
  wire       [1:0]    gateways_16_priority;
  reg                 gateways_16_ip;
  reg                 gateways_16_waitCompletion;
  wire                when_PlicGateway_l21_16;
  wire       [1:0]    gateways_17_priority;
  reg                 gateways_17_ip;
  reg                 gateways_17_waitCompletion;
  wire                when_PlicGateway_l21_17;
  wire       [1:0]    gateways_18_priority;
  reg                 gateways_18_ip;
  reg                 gateways_18_waitCompletion;
  wire                when_PlicGateway_l21_18;
  wire       [1:0]    gateways_19_priority;
  reg                 gateways_19_ip;
  reg                 gateways_19_waitCompletion;
  wire                when_PlicGateway_l21_19;
  wire       [1:0]    gateways_20_priority;
  reg                 gateways_20_ip;
  reg                 gateways_20_waitCompletion;
  wire                when_PlicGateway_l21_20;
  wire       [1:0]    gateways_21_priority;
  reg                 gateways_21_ip;
  reg                 gateways_21_waitCompletion;
  wire                when_PlicGateway_l21_21;
  wire       [1:0]    gateways_22_priority;
  reg                 gateways_22_ip;
  reg                 gateways_22_waitCompletion;
  wire                when_PlicGateway_l21_22;
  wire       [1:0]    gateways_23_priority;
  reg                 gateways_23_ip;
  reg                 gateways_23_waitCompletion;
  wire                when_PlicGateway_l21_23;
  wire       [1:0]    gateways_24_priority;
  reg                 gateways_24_ip;
  reg                 gateways_24_waitCompletion;
  wire                when_PlicGateway_l21_24;
  wire       [1:0]    gateways_25_priority;
  reg                 gateways_25_ip;
  reg                 gateways_25_waitCompletion;
  wire                when_PlicGateway_l21_25;
  wire       [1:0]    gateways_26_priority;
  reg                 gateways_26_ip;
  reg                 gateways_26_waitCompletion;
  wire                when_PlicGateway_l21_26;
  wire       [1:0]    gateways_27_priority;
  reg                 gateways_27_ip;
  reg                 gateways_27_waitCompletion;
  wire                when_PlicGateway_l21_27;
  wire       [1:0]    gateways_28_priority;
  reg                 gateways_28_ip;
  reg                 gateways_28_waitCompletion;
  wire                when_PlicGateway_l21_28;
  wire       [1:0]    gateways_29_priority;
  reg                 gateways_29_ip;
  reg                 gateways_29_waitCompletion;
  wire                when_PlicGateway_l21_29;
  wire       [1:0]    gateways_30_priority;
  reg                 gateways_30_ip;
  reg                 gateways_30_waitCompletion;
  wire                when_PlicGateway_l21_30;
  wire                targets_0_ie_0;
  wire                targets_0_ie_1;
  wire                targets_0_ie_2;
  wire                targets_0_ie_3;
  wire                targets_0_ie_4;
  wire                targets_0_ie_5;
  wire                targets_0_ie_6;
  wire                targets_0_ie_7;
  wire                targets_0_ie_8;
  wire                targets_0_ie_9;
  wire                targets_0_ie_10;
  wire                targets_0_ie_11;
  wire                targets_0_ie_12;
  wire                targets_0_ie_13;
  wire                targets_0_ie_14;
  wire                targets_0_ie_15;
  wire                targets_0_ie_16;
  wire                targets_0_ie_17;
  wire                targets_0_ie_18;
  wire                targets_0_ie_19;
  wire                targets_0_ie_20;
  wire                targets_0_ie_21;
  wire                targets_0_ie_22;
  wire                targets_0_ie_23;
  wire                targets_0_ie_24;
  wire                targets_0_ie_25;
  wire                targets_0_ie_26;
  wire                targets_0_ie_27;
  wire                targets_0_ie_28;
  wire                targets_0_ie_29;
  wire                targets_0_ie_30;
  wire       [1:0]    targets_0_threshold;
  wire       [1:0]    targets_0_requests_0_priority;
  wire       [4:0]    targets_0_requests_0_id;
  wire                targets_0_requests_0_valid;
  wire       [1:0]    targets_0_requests_1_priority;
  wire       [4:0]    targets_0_requests_1_id;
  wire                targets_0_requests_1_valid;
  wire       [1:0]    targets_0_requests_2_priority;
  wire       [4:0]    targets_0_requests_2_id;
  wire                targets_0_requests_2_valid;
  wire       [1:0]    targets_0_requests_3_priority;
  wire       [4:0]    targets_0_requests_3_id;
  wire                targets_0_requests_3_valid;
  wire       [1:0]    targets_0_requests_4_priority;
  wire       [4:0]    targets_0_requests_4_id;
  wire                targets_0_requests_4_valid;
  wire       [1:0]    targets_0_requests_5_priority;
  wire       [4:0]    targets_0_requests_5_id;
  wire                targets_0_requests_5_valid;
  wire       [1:0]    targets_0_requests_6_priority;
  wire       [4:0]    targets_0_requests_6_id;
  wire                targets_0_requests_6_valid;
  wire       [1:0]    targets_0_requests_7_priority;
  wire       [4:0]    targets_0_requests_7_id;
  wire                targets_0_requests_7_valid;
  wire       [1:0]    targets_0_requests_8_priority;
  wire       [4:0]    targets_0_requests_8_id;
  wire                targets_0_requests_8_valid;
  wire       [1:0]    targets_0_requests_9_priority;
  wire       [4:0]    targets_0_requests_9_id;
  wire                targets_0_requests_9_valid;
  wire       [1:0]    targets_0_requests_10_priority;
  wire       [4:0]    targets_0_requests_10_id;
  wire                targets_0_requests_10_valid;
  wire       [1:0]    targets_0_requests_11_priority;
  wire       [4:0]    targets_0_requests_11_id;
  wire                targets_0_requests_11_valid;
  wire       [1:0]    targets_0_requests_12_priority;
  wire       [4:0]    targets_0_requests_12_id;
  wire                targets_0_requests_12_valid;
  wire       [1:0]    targets_0_requests_13_priority;
  wire       [4:0]    targets_0_requests_13_id;
  wire                targets_0_requests_13_valid;
  wire       [1:0]    targets_0_requests_14_priority;
  wire       [4:0]    targets_0_requests_14_id;
  wire                targets_0_requests_14_valid;
  wire       [1:0]    targets_0_requests_15_priority;
  wire       [4:0]    targets_0_requests_15_id;
  wire                targets_0_requests_15_valid;
  wire       [1:0]    targets_0_requests_16_priority;
  wire       [4:0]    targets_0_requests_16_id;
  wire                targets_0_requests_16_valid;
  wire       [1:0]    targets_0_requests_17_priority;
  wire       [4:0]    targets_0_requests_17_id;
  wire                targets_0_requests_17_valid;
  wire       [1:0]    targets_0_requests_18_priority;
  wire       [4:0]    targets_0_requests_18_id;
  wire                targets_0_requests_18_valid;
  wire       [1:0]    targets_0_requests_19_priority;
  wire       [4:0]    targets_0_requests_19_id;
  wire                targets_0_requests_19_valid;
  wire       [1:0]    targets_0_requests_20_priority;
  wire       [4:0]    targets_0_requests_20_id;
  wire                targets_0_requests_20_valid;
  wire       [1:0]    targets_0_requests_21_priority;
  wire       [4:0]    targets_0_requests_21_id;
  wire                targets_0_requests_21_valid;
  wire       [1:0]    targets_0_requests_22_priority;
  wire       [4:0]    targets_0_requests_22_id;
  wire                targets_0_requests_22_valid;
  wire       [1:0]    targets_0_requests_23_priority;
  wire       [4:0]    targets_0_requests_23_id;
  wire                targets_0_requests_23_valid;
  wire       [1:0]    targets_0_requests_24_priority;
  wire       [4:0]    targets_0_requests_24_id;
  wire                targets_0_requests_24_valid;
  wire       [1:0]    targets_0_requests_25_priority;
  wire       [4:0]    targets_0_requests_25_id;
  wire                targets_0_requests_25_valid;
  wire       [1:0]    targets_0_requests_26_priority;
  wire       [4:0]    targets_0_requests_26_id;
  wire                targets_0_requests_26_valid;
  wire       [1:0]    targets_0_requests_27_priority;
  wire       [4:0]    targets_0_requests_27_id;
  wire                targets_0_requests_27_valid;
  wire       [1:0]    targets_0_requests_28_priority;
  wire       [4:0]    targets_0_requests_28_id;
  wire                targets_0_requests_28_valid;
  wire       [1:0]    targets_0_requests_29_priority;
  wire       [4:0]    targets_0_requests_29_id;
  wire                targets_0_requests_29_valid;
  wire       [1:0]    targets_0_requests_30_priority;
  wire       [4:0]    targets_0_requests_30_id;
  wire                targets_0_requests_30_valid;
  wire       [1:0]    targets_0_requests_31_priority;
  wire       [4:0]    targets_0_requests_31_id;
  wire                targets_0_requests_31_valid;
  wire                _zz_targets_0_bestRequest_id;
  wire       [1:0]    _zz_targets_0_bestRequest_id_1;
  wire                _zz_targets_0_bestRequest_id_2;
  wire                _zz_targets_0_bestRequest_id_3;
  wire       [1:0]    _zz_targets_0_bestRequest_id_4;
  wire                _zz_targets_0_bestRequest_id_5;
  wire                _zz_targets_0_bestRequest_id_6;
  wire       [1:0]    _zz_targets_0_bestRequest_id_7;
  wire                _zz_targets_0_bestRequest_id_8;
  wire                _zz_targets_0_bestRequest_id_9;
  wire       [1:0]    _zz_targets_0_bestRequest_id_10;
  wire                _zz_targets_0_bestRequest_id_11;
  wire                _zz_targets_0_bestRequest_id_12;
  wire       [1:0]    _zz_targets_0_bestRequest_id_13;
  wire                _zz_targets_0_bestRequest_id_14;
  wire                _zz_targets_0_bestRequest_id_15;
  wire       [1:0]    _zz_targets_0_bestRequest_id_16;
  wire                _zz_targets_0_bestRequest_id_17;
  wire                _zz_targets_0_bestRequest_id_18;
  wire       [1:0]    _zz_targets_0_bestRequest_id_19;
  wire                _zz_targets_0_bestRequest_id_20;
  wire                _zz_targets_0_bestRequest_id_21;
  wire       [1:0]    _zz_targets_0_bestRequest_id_22;
  wire                _zz_targets_0_bestRequest_id_23;
  wire                _zz_targets_0_bestRequest_id_24;
  wire       [1:0]    _zz_targets_0_bestRequest_id_25;
  wire                _zz_targets_0_bestRequest_id_26;
  wire                _zz_targets_0_bestRequest_id_27;
  wire       [1:0]    _zz_targets_0_bestRequest_id_28;
  wire                _zz_targets_0_bestRequest_id_29;
  wire                _zz_targets_0_bestRequest_id_30;
  wire       [1:0]    _zz_targets_0_bestRequest_id_31;
  wire                _zz_targets_0_bestRequest_id_32;
  wire                _zz_targets_0_bestRequest_id_33;
  wire       [1:0]    _zz_targets_0_bestRequest_id_34;
  wire                _zz_targets_0_bestRequest_id_35;
  wire                _zz_targets_0_bestRequest_id_36;
  wire       [1:0]    _zz_targets_0_bestRequest_id_37;
  wire                _zz_targets_0_bestRequest_id_38;
  wire                _zz_targets_0_bestRequest_id_39;
  wire       [1:0]    _zz_targets_0_bestRequest_id_40;
  wire                _zz_targets_0_bestRequest_id_41;
  wire                _zz_targets_0_bestRequest_id_42;
  wire       [1:0]    _zz_targets_0_bestRequest_id_43;
  wire                _zz_targets_0_bestRequest_id_44;
  wire                _zz_targets_0_bestRequest_id_45;
  wire       [1:0]    _zz_targets_0_bestRequest_id_46;
  wire                _zz_targets_0_bestRequest_id_47;
  wire                _zz_targets_0_bestRequest_id_48;
  wire       [1:0]    _zz_targets_0_bestRequest_id_49;
  wire                _zz_targets_0_bestRequest_id_50;
  wire                _zz_targets_0_bestRequest_id_51;
  wire       [1:0]    _zz_targets_0_bestRequest_id_52;
  wire                _zz_targets_0_bestRequest_id_53;
  wire                _zz_targets_0_bestRequest_id_54;
  wire       [1:0]    _zz_targets_0_bestRequest_id_55;
  wire                _zz_targets_0_bestRequest_id_56;
  wire                _zz_targets_0_bestRequest_id_57;
  wire       [1:0]    _zz_targets_0_bestRequest_id_58;
  wire                _zz_targets_0_bestRequest_id_59;
  wire                _zz_targets_0_bestRequest_id_60;
  wire       [1:0]    _zz_targets_0_bestRequest_id_61;
  wire                _zz_targets_0_bestRequest_id_62;
  wire                _zz_targets_0_bestRequest_id_63;
  wire       [1:0]    _zz_targets_0_bestRequest_id_64;
  wire                _zz_targets_0_bestRequest_id_65;
  wire                _zz_targets_0_bestRequest_id_66;
  wire       [1:0]    _zz_targets_0_bestRequest_id_67;
  wire                _zz_targets_0_bestRequest_id_68;
  wire                _zz_targets_0_bestRequest_id_69;
  wire       [1:0]    _zz_targets_0_bestRequest_id_70;
  wire                _zz_targets_0_bestRequest_id_71;
  wire                _zz_targets_0_bestRequest_id_72;
  wire       [1:0]    _zz_targets_0_bestRequest_priority;
  wire                _zz_targets_0_bestRequest_id_73;
  wire                _zz_targets_0_bestRequest_id_74;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_1;
  wire                _zz_targets_0_bestRequest_id_75;
  wire                _zz_targets_0_bestRequest_id_76;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_2;
  wire                _zz_targets_0_bestRequest_id_77;
  wire                _zz_targets_0_bestRequest_id_78;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_3;
  wire                _zz_targets_0_bestRequest_id_79;
  wire                _zz_targets_0_bestRequest_id_80;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_4;
  wire                _zz_targets_0_bestRequest_valid;
  wire                _zz_targets_0_bestRequest_id_81;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_5;
  wire                _zz_targets_0_bestRequest_valid_1;
  wire                _zz_targets_0_bestRequest_priority_6;
  reg        [1:0]    targets_0_bestRequest_priority;
  reg        [4:0]    targets_0_bestRequest_id;
  reg                 targets_0_bestRequest_valid;
  wire                targets_0_iep;
  wire       [4:0]    targets_0_claim;
  wire                targets_1_ie_0;
  wire                targets_1_ie_1;
  wire                targets_1_ie_2;
  wire                targets_1_ie_3;
  wire                targets_1_ie_4;
  wire                targets_1_ie_5;
  wire                targets_1_ie_6;
  wire                targets_1_ie_7;
  wire                targets_1_ie_8;
  wire                targets_1_ie_9;
  wire                targets_1_ie_10;
  wire                targets_1_ie_11;
  wire                targets_1_ie_12;
  wire                targets_1_ie_13;
  wire                targets_1_ie_14;
  wire                targets_1_ie_15;
  wire                targets_1_ie_16;
  wire                targets_1_ie_17;
  wire                targets_1_ie_18;
  wire                targets_1_ie_19;
  wire                targets_1_ie_20;
  wire                targets_1_ie_21;
  wire                targets_1_ie_22;
  wire                targets_1_ie_23;
  wire                targets_1_ie_24;
  wire                targets_1_ie_25;
  wire                targets_1_ie_26;
  wire                targets_1_ie_27;
  wire                targets_1_ie_28;
  wire                targets_1_ie_29;
  wire                targets_1_ie_30;
  wire       [1:0]    targets_1_threshold;
  wire       [1:0]    targets_1_requests_0_priority;
  wire       [4:0]    targets_1_requests_0_id;
  wire                targets_1_requests_0_valid;
  wire       [1:0]    targets_1_requests_1_priority;
  wire       [4:0]    targets_1_requests_1_id;
  wire                targets_1_requests_1_valid;
  wire       [1:0]    targets_1_requests_2_priority;
  wire       [4:0]    targets_1_requests_2_id;
  wire                targets_1_requests_2_valid;
  wire       [1:0]    targets_1_requests_3_priority;
  wire       [4:0]    targets_1_requests_3_id;
  wire                targets_1_requests_3_valid;
  wire       [1:0]    targets_1_requests_4_priority;
  wire       [4:0]    targets_1_requests_4_id;
  wire                targets_1_requests_4_valid;
  wire       [1:0]    targets_1_requests_5_priority;
  wire       [4:0]    targets_1_requests_5_id;
  wire                targets_1_requests_5_valid;
  wire       [1:0]    targets_1_requests_6_priority;
  wire       [4:0]    targets_1_requests_6_id;
  wire                targets_1_requests_6_valid;
  wire       [1:0]    targets_1_requests_7_priority;
  wire       [4:0]    targets_1_requests_7_id;
  wire                targets_1_requests_7_valid;
  wire       [1:0]    targets_1_requests_8_priority;
  wire       [4:0]    targets_1_requests_8_id;
  wire                targets_1_requests_8_valid;
  wire       [1:0]    targets_1_requests_9_priority;
  wire       [4:0]    targets_1_requests_9_id;
  wire                targets_1_requests_9_valid;
  wire       [1:0]    targets_1_requests_10_priority;
  wire       [4:0]    targets_1_requests_10_id;
  wire                targets_1_requests_10_valid;
  wire       [1:0]    targets_1_requests_11_priority;
  wire       [4:0]    targets_1_requests_11_id;
  wire                targets_1_requests_11_valid;
  wire       [1:0]    targets_1_requests_12_priority;
  wire       [4:0]    targets_1_requests_12_id;
  wire                targets_1_requests_12_valid;
  wire       [1:0]    targets_1_requests_13_priority;
  wire       [4:0]    targets_1_requests_13_id;
  wire                targets_1_requests_13_valid;
  wire       [1:0]    targets_1_requests_14_priority;
  wire       [4:0]    targets_1_requests_14_id;
  wire                targets_1_requests_14_valid;
  wire       [1:0]    targets_1_requests_15_priority;
  wire       [4:0]    targets_1_requests_15_id;
  wire                targets_1_requests_15_valid;
  wire       [1:0]    targets_1_requests_16_priority;
  wire       [4:0]    targets_1_requests_16_id;
  wire                targets_1_requests_16_valid;
  wire       [1:0]    targets_1_requests_17_priority;
  wire       [4:0]    targets_1_requests_17_id;
  wire                targets_1_requests_17_valid;
  wire       [1:0]    targets_1_requests_18_priority;
  wire       [4:0]    targets_1_requests_18_id;
  wire                targets_1_requests_18_valid;
  wire       [1:0]    targets_1_requests_19_priority;
  wire       [4:0]    targets_1_requests_19_id;
  wire                targets_1_requests_19_valid;
  wire       [1:0]    targets_1_requests_20_priority;
  wire       [4:0]    targets_1_requests_20_id;
  wire                targets_1_requests_20_valid;
  wire       [1:0]    targets_1_requests_21_priority;
  wire       [4:0]    targets_1_requests_21_id;
  wire                targets_1_requests_21_valid;
  wire       [1:0]    targets_1_requests_22_priority;
  wire       [4:0]    targets_1_requests_22_id;
  wire                targets_1_requests_22_valid;
  wire       [1:0]    targets_1_requests_23_priority;
  wire       [4:0]    targets_1_requests_23_id;
  wire                targets_1_requests_23_valid;
  wire       [1:0]    targets_1_requests_24_priority;
  wire       [4:0]    targets_1_requests_24_id;
  wire                targets_1_requests_24_valid;
  wire       [1:0]    targets_1_requests_25_priority;
  wire       [4:0]    targets_1_requests_25_id;
  wire                targets_1_requests_25_valid;
  wire       [1:0]    targets_1_requests_26_priority;
  wire       [4:0]    targets_1_requests_26_id;
  wire                targets_1_requests_26_valid;
  wire       [1:0]    targets_1_requests_27_priority;
  wire       [4:0]    targets_1_requests_27_id;
  wire                targets_1_requests_27_valid;
  wire       [1:0]    targets_1_requests_28_priority;
  wire       [4:0]    targets_1_requests_28_id;
  wire                targets_1_requests_28_valid;
  wire       [1:0]    targets_1_requests_29_priority;
  wire       [4:0]    targets_1_requests_29_id;
  wire                targets_1_requests_29_valid;
  wire       [1:0]    targets_1_requests_30_priority;
  wire       [4:0]    targets_1_requests_30_id;
  wire                targets_1_requests_30_valid;
  wire       [1:0]    targets_1_requests_31_priority;
  wire       [4:0]    targets_1_requests_31_id;
  wire                targets_1_requests_31_valid;
  wire                _zz_targets_1_bestRequest_id;
  wire       [1:0]    _zz_targets_1_bestRequest_id_1;
  wire                _zz_targets_1_bestRequest_id_2;
  wire                _zz_targets_1_bestRequest_id_3;
  wire       [1:0]    _zz_targets_1_bestRequest_id_4;
  wire                _zz_targets_1_bestRequest_id_5;
  wire                _zz_targets_1_bestRequest_id_6;
  wire       [1:0]    _zz_targets_1_bestRequest_id_7;
  wire                _zz_targets_1_bestRequest_id_8;
  wire                _zz_targets_1_bestRequest_id_9;
  wire       [1:0]    _zz_targets_1_bestRequest_id_10;
  wire                _zz_targets_1_bestRequest_id_11;
  wire                _zz_targets_1_bestRequest_id_12;
  wire       [1:0]    _zz_targets_1_bestRequest_id_13;
  wire                _zz_targets_1_bestRequest_id_14;
  wire                _zz_targets_1_bestRequest_id_15;
  wire       [1:0]    _zz_targets_1_bestRequest_id_16;
  wire                _zz_targets_1_bestRequest_id_17;
  wire                _zz_targets_1_bestRequest_id_18;
  wire       [1:0]    _zz_targets_1_bestRequest_id_19;
  wire                _zz_targets_1_bestRequest_id_20;
  wire                _zz_targets_1_bestRequest_id_21;
  wire       [1:0]    _zz_targets_1_bestRequest_id_22;
  wire                _zz_targets_1_bestRequest_id_23;
  wire                _zz_targets_1_bestRequest_id_24;
  wire       [1:0]    _zz_targets_1_bestRequest_id_25;
  wire                _zz_targets_1_bestRequest_id_26;
  wire                _zz_targets_1_bestRequest_id_27;
  wire       [1:0]    _zz_targets_1_bestRequest_id_28;
  wire                _zz_targets_1_bestRequest_id_29;
  wire                _zz_targets_1_bestRequest_id_30;
  wire       [1:0]    _zz_targets_1_bestRequest_id_31;
  wire                _zz_targets_1_bestRequest_id_32;
  wire                _zz_targets_1_bestRequest_id_33;
  wire       [1:0]    _zz_targets_1_bestRequest_id_34;
  wire                _zz_targets_1_bestRequest_id_35;
  wire                _zz_targets_1_bestRequest_id_36;
  wire       [1:0]    _zz_targets_1_bestRequest_id_37;
  wire                _zz_targets_1_bestRequest_id_38;
  wire                _zz_targets_1_bestRequest_id_39;
  wire       [1:0]    _zz_targets_1_bestRequest_id_40;
  wire                _zz_targets_1_bestRequest_id_41;
  wire                _zz_targets_1_bestRequest_id_42;
  wire       [1:0]    _zz_targets_1_bestRequest_id_43;
  wire                _zz_targets_1_bestRequest_id_44;
  wire                _zz_targets_1_bestRequest_id_45;
  wire       [1:0]    _zz_targets_1_bestRequest_id_46;
  wire                _zz_targets_1_bestRequest_id_47;
  wire                _zz_targets_1_bestRequest_id_48;
  wire       [1:0]    _zz_targets_1_bestRequest_id_49;
  wire                _zz_targets_1_bestRequest_id_50;
  wire                _zz_targets_1_bestRequest_id_51;
  wire       [1:0]    _zz_targets_1_bestRequest_id_52;
  wire                _zz_targets_1_bestRequest_id_53;
  wire                _zz_targets_1_bestRequest_id_54;
  wire       [1:0]    _zz_targets_1_bestRequest_id_55;
  wire                _zz_targets_1_bestRequest_id_56;
  wire                _zz_targets_1_bestRequest_id_57;
  wire       [1:0]    _zz_targets_1_bestRequest_id_58;
  wire                _zz_targets_1_bestRequest_id_59;
  wire                _zz_targets_1_bestRequest_id_60;
  wire       [1:0]    _zz_targets_1_bestRequest_id_61;
  wire                _zz_targets_1_bestRequest_id_62;
  wire                _zz_targets_1_bestRequest_id_63;
  wire       [1:0]    _zz_targets_1_bestRequest_id_64;
  wire                _zz_targets_1_bestRequest_id_65;
  wire                _zz_targets_1_bestRequest_id_66;
  wire       [1:0]    _zz_targets_1_bestRequest_id_67;
  wire                _zz_targets_1_bestRequest_id_68;
  wire                _zz_targets_1_bestRequest_id_69;
  wire       [1:0]    _zz_targets_1_bestRequest_id_70;
  wire                _zz_targets_1_bestRequest_id_71;
  wire                _zz_targets_1_bestRequest_id_72;
  wire       [1:0]    _zz_targets_1_bestRequest_priority;
  wire                _zz_targets_1_bestRequest_id_73;
  wire                _zz_targets_1_bestRequest_id_74;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_1;
  wire                _zz_targets_1_bestRequest_id_75;
  wire                _zz_targets_1_bestRequest_id_76;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_2;
  wire                _zz_targets_1_bestRequest_id_77;
  wire                _zz_targets_1_bestRequest_id_78;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_3;
  wire                _zz_targets_1_bestRequest_id_79;
  wire                _zz_targets_1_bestRequest_id_80;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_4;
  wire                _zz_targets_1_bestRequest_valid;
  wire                _zz_targets_1_bestRequest_id_81;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_5;
  wire                _zz_targets_1_bestRequest_valid_1;
  wire                _zz_targets_1_bestRequest_priority_6;
  reg        [1:0]    targets_1_bestRequest_priority;
  reg        [4:0]    targets_1_bestRequest_id;
  reg                 targets_1_bestRequest_valid;
  wire                targets_1_iep;
  wire       [4:0]    targets_1_claim;
  wire                bus_readErrorFlag;
  wire                bus_writeErrorFlag;
  reg                 bus_readHaltRequest;
  wire                bus_writeHaltRequest;
  wire                bus_writeJoinEvent_valid;
  wire                bus_writeJoinEvent_ready;
  wire                bus_writeOccur;
  reg        [1:0]    bus_writeRsp_resp;
  wire                bus_writeJoinEvent_translated_valid;
  wire                bus_writeJoinEvent_translated_ready;
  wire       [1:0]    bus_writeJoinEvent_translated_payload_resp;
  wire                _zz_bus_writeJoinEvent_translated_ready;
  wire                _zz_bus_writeJoinEvent_translated_ready_1;
  wire                _zz_io_bus_b_valid;
  reg                 _zz_io_bus_b_valid_1;
  reg        [1:0]    _zz_io_bus_b_payload_resp;
  wire                bus_readDataStage_valid;
  wire                bus_readDataStage_ready;
  wire       [21:0]   bus_readDataStage_payload_addr;
  wire       [2:0]    bus_readDataStage_payload_prot;
  reg                 io_bus_ar_rValid;
  wire                bus_readDataStage_fire;
  reg        [21:0]   io_bus_ar_rData_addr;
  reg        [2:0]    io_bus_ar_rData_prot;
  reg        [31:0]   bus_readRsp_data;
  reg        [1:0]    bus_readRsp_resp;
  wire                _zz_io_bus_r_valid;
  wire       [21:0]   bus_readAddressMasked;
  wire       [21:0]   bus_writeAddressMasked;
  wire                bus_readOccur;
  reg        [1:0]    _zz_gateways_0_priority;
  reg        [1:0]    _zz_gateways_1_priority;
  reg        [1:0]    _zz_gateways_2_priority;
  reg        [1:0]    _zz_gateways_3_priority;
  reg        [1:0]    _zz_gateways_4_priority;
  reg        [1:0]    _zz_gateways_5_priority;
  reg        [1:0]    _zz_gateways_6_priority;
  reg        [1:0]    _zz_gateways_7_priority;
  reg        [1:0]    _zz_gateways_8_priority;
  reg        [1:0]    _zz_gateways_9_priority;
  reg        [1:0]    _zz_gateways_10_priority;
  reg        [1:0]    _zz_gateways_11_priority;
  reg        [1:0]    _zz_gateways_12_priority;
  reg        [1:0]    _zz_gateways_13_priority;
  reg        [1:0]    _zz_gateways_14_priority;
  reg        [1:0]    _zz_gateways_15_priority;
  reg        [1:0]    _zz_gateways_16_priority;
  reg        [1:0]    _zz_gateways_17_priority;
  reg        [1:0]    _zz_gateways_18_priority;
  reg        [1:0]    _zz_gateways_19_priority;
  reg        [1:0]    _zz_gateways_20_priority;
  reg        [1:0]    _zz_gateways_21_priority;
  reg        [1:0]    _zz_gateways_22_priority;
  reg        [1:0]    _zz_gateways_23_priority;
  reg        [1:0]    _zz_gateways_24_priority;
  reg        [1:0]    _zz_gateways_25_priority;
  reg        [1:0]    _zz_gateways_26_priority;
  reg        [1:0]    _zz_gateways_27_priority;
  reg        [1:0]    _zz_gateways_28_priority;
  reg        [1:0]    _zz_gateways_29_priority;
  reg        [1:0]    _zz_gateways_30_priority;
  reg                 mapping_claim_valid;
  reg        [4:0]    mapping_claim_payload;
  reg                 mapping_completion_valid;
  reg        [4:0]    mapping_completion_payload;
  reg                 mapping_coherencyStall_willIncrement;
  wire                mapping_coherencyStall_willClear;
  reg        [0:0]    mapping_coherencyStall_valueNext;
  reg        [0:0]    mapping_coherencyStall_value;
  wire                mapping_coherencyStall_willOverflowIfInc;
  wire                mapping_coherencyStall_willOverflow;
  wire                when_PlicMapper_l122;
  reg        [1:0]    _zz_targets_0_threshold;
  reg                 mapping_targetMapping_0_targetCompletion_valid;
  wire       [4:0]    mapping_targetMapping_0_targetCompletion_payload;
  reg                 _zz_targets_0_ie_0;
  reg                 _zz_targets_0_ie_1;
  reg                 _zz_targets_0_ie_2;
  reg                 _zz_targets_0_ie_3;
  reg                 _zz_targets_0_ie_4;
  reg                 _zz_targets_0_ie_5;
  reg                 _zz_targets_0_ie_6;
  reg                 _zz_targets_0_ie_7;
  reg                 _zz_targets_0_ie_8;
  reg                 _zz_targets_0_ie_9;
  reg                 _zz_targets_0_ie_10;
  reg                 _zz_targets_0_ie_11;
  reg                 _zz_targets_0_ie_12;
  reg                 _zz_targets_0_ie_13;
  reg                 _zz_targets_0_ie_14;
  reg                 _zz_targets_0_ie_15;
  reg                 _zz_targets_0_ie_16;
  reg                 _zz_targets_0_ie_17;
  reg                 _zz_targets_0_ie_18;
  reg                 _zz_targets_0_ie_19;
  reg                 _zz_targets_0_ie_20;
  reg                 _zz_targets_0_ie_21;
  reg                 _zz_targets_0_ie_22;
  reg                 _zz_targets_0_ie_23;
  reg                 _zz_targets_0_ie_24;
  reg                 _zz_targets_0_ie_25;
  reg                 _zz_targets_0_ie_26;
  reg                 _zz_targets_0_ie_27;
  reg                 _zz_targets_0_ie_28;
  reg                 _zz_targets_0_ie_29;
  reg                 _zz_targets_0_ie_30;
  reg        [1:0]    _zz_targets_1_threshold;
  reg                 mapping_targetMapping_1_targetCompletion_valid;
  wire       [4:0]    mapping_targetMapping_1_targetCompletion_payload;
  reg                 _zz_targets_1_ie_0;
  reg                 _zz_targets_1_ie_1;
  reg                 _zz_targets_1_ie_2;
  reg                 _zz_targets_1_ie_3;
  reg                 _zz_targets_1_ie_4;
  reg                 _zz_targets_1_ie_5;
  reg                 _zz_targets_1_ie_6;
  reg                 _zz_targets_1_ie_7;
  reg                 _zz_targets_1_ie_8;
  reg                 _zz_targets_1_ie_9;
  reg                 _zz_targets_1_ie_10;
  reg                 _zz_targets_1_ie_11;
  reg                 _zz_targets_1_ie_12;
  reg                 _zz_targets_1_ie_13;
  reg                 _zz_targets_1_ie_14;
  reg                 _zz_targets_1_ie_15;
  reg                 _zz_targets_1_ie_16;
  reg                 _zz_targets_1_ie_17;
  reg                 _zz_targets_1_ie_18;
  reg                 _zz_targets_1_ie_19;
  reg                 _zz_targets_1_ie_20;
  reg                 _zz_targets_1_ie_21;
  reg                 _zz_targets_1_ie_22;
  reg                 _zz_targets_1_ie_23;
  reg                 _zz_targets_1_ie_24;
  reg                 _zz_targets_1_ie_25;
  reg                 _zz_targets_1_ie_26;
  reg                 _zz_targets_1_ie_27;
  reg                 _zz_targets_1_ie_28;
  reg                 _zz_targets_1_ie_29;
  reg                 _zz_targets_1_ie_30;
  wire                when_AxiLite4SlaveFactory_l68;
  wire                when_AxiLite4SlaveFactory_l86;

  assign _zz_targets_0_bestRequest_id_82 = (_zz_targets_0_bestRequest_id ? targets_0_requests_0_id : targets_0_requests_1_id);
  assign _zz_targets_0_bestRequest_id_83 = (_zz_targets_0_bestRequest_id_3 ? targets_0_requests_2_id : targets_0_requests_3_id);
  assign _zz_targets_0_bestRequest_id_84 = (_zz_targets_0_bestRequest_id_6 ? targets_0_requests_4_id : targets_0_requests_5_id);
  assign _zz_targets_0_bestRequest_id_85 = (_zz_targets_0_bestRequest_id_9 ? targets_0_requests_6_id : targets_0_requests_7_id);
  assign _zz_targets_0_bestRequest_id_86 = (_zz_targets_0_bestRequest_id_12 ? targets_0_requests_8_id : targets_0_requests_9_id);
  assign _zz_targets_0_bestRequest_id_87 = (_zz_targets_0_bestRequest_id_15 ? targets_0_requests_10_id : targets_0_requests_11_id);
  assign _zz_targets_0_bestRequest_id_88 = (_zz_targets_0_bestRequest_id_18 ? targets_0_requests_12_id : targets_0_requests_13_id);
  assign _zz_targets_0_bestRequest_id_89 = (_zz_targets_0_bestRequest_id_21 ? targets_0_requests_14_id : targets_0_requests_15_id);
  assign _zz_targets_0_bestRequest_id_90 = (_zz_targets_0_bestRequest_id_24 ? targets_0_requests_16_id : targets_0_requests_17_id);
  assign _zz_targets_0_bestRequest_id_91 = (_zz_targets_0_bestRequest_id_27 ? targets_0_requests_18_id : targets_0_requests_19_id);
  assign _zz_targets_0_bestRequest_id_92 = (_zz_targets_0_bestRequest_id_30 ? targets_0_requests_20_id : targets_0_requests_21_id);
  assign _zz_targets_0_bestRequest_id_93 = (_zz_targets_0_bestRequest_id_33 ? targets_0_requests_22_id : targets_0_requests_23_id);
  assign _zz_targets_0_bestRequest_id_94 = (_zz_targets_0_bestRequest_id_36 ? targets_0_requests_24_id : targets_0_requests_25_id);
  assign _zz_targets_0_bestRequest_id_95 = (_zz_targets_0_bestRequest_id_39 ? targets_0_requests_26_id : targets_0_requests_27_id);
  assign _zz_targets_0_bestRequest_id_96 = (_zz_targets_0_bestRequest_id_42 ? targets_0_requests_28_id : targets_0_requests_29_id);
  assign _zz_targets_0_bestRequest_id_97 = (_zz_targets_0_bestRequest_id_45 ? targets_0_requests_30_id : targets_0_requests_31_id);
  assign _zz_targets_1_bestRequest_id_82 = (_zz_targets_1_bestRequest_id ? targets_1_requests_0_id : targets_1_requests_1_id);
  assign _zz_targets_1_bestRequest_id_83 = (_zz_targets_1_bestRequest_id_3 ? targets_1_requests_2_id : targets_1_requests_3_id);
  assign _zz_targets_1_bestRequest_id_84 = (_zz_targets_1_bestRequest_id_6 ? targets_1_requests_4_id : targets_1_requests_5_id);
  assign _zz_targets_1_bestRequest_id_85 = (_zz_targets_1_bestRequest_id_9 ? targets_1_requests_6_id : targets_1_requests_7_id);
  assign _zz_targets_1_bestRequest_id_86 = (_zz_targets_1_bestRequest_id_12 ? targets_1_requests_8_id : targets_1_requests_9_id);
  assign _zz_targets_1_bestRequest_id_87 = (_zz_targets_1_bestRequest_id_15 ? targets_1_requests_10_id : targets_1_requests_11_id);
  assign _zz_targets_1_bestRequest_id_88 = (_zz_targets_1_bestRequest_id_18 ? targets_1_requests_12_id : targets_1_requests_13_id);
  assign _zz_targets_1_bestRequest_id_89 = (_zz_targets_1_bestRequest_id_21 ? targets_1_requests_14_id : targets_1_requests_15_id);
  assign _zz_targets_1_bestRequest_id_90 = (_zz_targets_1_bestRequest_id_24 ? targets_1_requests_16_id : targets_1_requests_17_id);
  assign _zz_targets_1_bestRequest_id_91 = (_zz_targets_1_bestRequest_id_27 ? targets_1_requests_18_id : targets_1_requests_19_id);
  assign _zz_targets_1_bestRequest_id_92 = (_zz_targets_1_bestRequest_id_30 ? targets_1_requests_20_id : targets_1_requests_21_id);
  assign _zz_targets_1_bestRequest_id_93 = (_zz_targets_1_bestRequest_id_33 ? targets_1_requests_22_id : targets_1_requests_23_id);
  assign _zz_targets_1_bestRequest_id_94 = (_zz_targets_1_bestRequest_id_36 ? targets_1_requests_24_id : targets_1_requests_25_id);
  assign _zz_targets_1_bestRequest_id_95 = (_zz_targets_1_bestRequest_id_39 ? targets_1_requests_26_id : targets_1_requests_27_id);
  assign _zz_targets_1_bestRequest_id_96 = (_zz_targets_1_bestRequest_id_42 ? targets_1_requests_28_id : targets_1_requests_29_id);
  assign _zz_targets_1_bestRequest_id_97 = (_zz_targets_1_bestRequest_id_45 ? targets_1_requests_30_id : targets_1_requests_31_id);
  assign _zz_gateways_0_ip = io_sources[0];
  assign _zz_gateways_1_ip = io_sources[1];
  assign _zz_gateways_2_ip = io_sources[2];
  assign _zz_gateways_3_ip = io_sources[3];
  assign _zz_gateways_4_ip = io_sources[4];
  assign _zz_gateways_5_ip = io_sources[5];
  assign _zz_gateways_6_ip = io_sources[6];
  assign _zz_gateways_7_ip = io_sources[7];
  assign _zz_gateways_8_ip = io_sources[8];
  assign _zz_gateways_9_ip = io_sources[9];
  assign _zz_gateways_10_ip = io_sources[10];
  assign _zz_gateways_11_ip = io_sources[11];
  assign _zz_gateways_12_ip = io_sources[12];
  assign _zz_gateways_13_ip = io_sources[13];
  assign _zz_gateways_14_ip = io_sources[14];
  assign _zz_gateways_15_ip = io_sources[15];
  assign _zz_gateways_16_ip = io_sources[16];
  assign _zz_gateways_17_ip = io_sources[17];
  assign _zz_gateways_18_ip = io_sources[18];
  assign _zz_gateways_19_ip = io_sources[19];
  assign _zz_gateways_20_ip = io_sources[20];
  assign _zz_gateways_21_ip = io_sources[21];
  assign _zz_gateways_22_ip = io_sources[22];
  assign _zz_gateways_23_ip = io_sources[23];
  assign _zz_gateways_24_ip = io_sources[24];
  assign _zz_gateways_25_ip = io_sources[25];
  assign _zz_gateways_26_ip = io_sources[26];
  assign _zz_gateways_27_ip = io_sources[27];
  assign _zz_gateways_28_ip = io_sources[28];
  assign _zz_gateways_29_ip = io_sources[29];
  assign _zz_gateways_30_ip = io_sources[30];
  assign when_PlicGateway_l21 = (! gateways_0_waitCompletion);
  assign when_PlicGateway_l21_1 = (! gateways_1_waitCompletion);
  assign when_PlicGateway_l21_2 = (! gateways_2_waitCompletion);
  assign when_PlicGateway_l21_3 = (! gateways_3_waitCompletion);
  assign when_PlicGateway_l21_4 = (! gateways_4_waitCompletion);
  assign when_PlicGateway_l21_5 = (! gateways_5_waitCompletion);
  assign when_PlicGateway_l21_6 = (! gateways_6_waitCompletion);
  assign when_PlicGateway_l21_7 = (! gateways_7_waitCompletion);
  assign when_PlicGateway_l21_8 = (! gateways_8_waitCompletion);
  assign when_PlicGateway_l21_9 = (! gateways_9_waitCompletion);
  assign when_PlicGateway_l21_10 = (! gateways_10_waitCompletion);
  assign when_PlicGateway_l21_11 = (! gateways_11_waitCompletion);
  assign when_PlicGateway_l21_12 = (! gateways_12_waitCompletion);
  assign when_PlicGateway_l21_13 = (! gateways_13_waitCompletion);
  assign when_PlicGateway_l21_14 = (! gateways_14_waitCompletion);
  assign when_PlicGateway_l21_15 = (! gateways_15_waitCompletion);
  assign when_PlicGateway_l21_16 = (! gateways_16_waitCompletion);
  assign when_PlicGateway_l21_17 = (! gateways_17_waitCompletion);
  assign when_PlicGateway_l21_18 = (! gateways_18_waitCompletion);
  assign when_PlicGateway_l21_19 = (! gateways_19_waitCompletion);
  assign when_PlicGateway_l21_20 = (! gateways_20_waitCompletion);
  assign when_PlicGateway_l21_21 = (! gateways_21_waitCompletion);
  assign when_PlicGateway_l21_22 = (! gateways_22_waitCompletion);
  assign when_PlicGateway_l21_23 = (! gateways_23_waitCompletion);
  assign when_PlicGateway_l21_24 = (! gateways_24_waitCompletion);
  assign when_PlicGateway_l21_25 = (! gateways_25_waitCompletion);
  assign when_PlicGateway_l21_26 = (! gateways_26_waitCompletion);
  assign when_PlicGateway_l21_27 = (! gateways_27_waitCompletion);
  assign when_PlicGateway_l21_28 = (! gateways_28_waitCompletion);
  assign when_PlicGateway_l21_29 = (! gateways_29_waitCompletion);
  assign when_PlicGateway_l21_30 = (! gateways_30_waitCompletion);
  assign targets_0_requests_0_priority = 2'b00;
  assign targets_0_requests_0_id = 5'h00;
  assign targets_0_requests_0_valid = 1'b1;
  assign targets_0_requests_1_priority = gateways_0_priority;
  assign targets_0_requests_1_id = 5'h01;
  assign targets_0_requests_1_valid = (gateways_0_ip && targets_0_ie_0);
  assign targets_0_requests_2_priority = gateways_1_priority;
  assign targets_0_requests_2_id = 5'h02;
  assign targets_0_requests_2_valid = (gateways_1_ip && targets_0_ie_1);
  assign targets_0_requests_3_priority = gateways_2_priority;
  assign targets_0_requests_3_id = 5'h03;
  assign targets_0_requests_3_valid = (gateways_2_ip && targets_0_ie_2);
  assign targets_0_requests_4_priority = gateways_3_priority;
  assign targets_0_requests_4_id = 5'h04;
  assign targets_0_requests_4_valid = (gateways_3_ip && targets_0_ie_3);
  assign targets_0_requests_5_priority = gateways_4_priority;
  assign targets_0_requests_5_id = 5'h05;
  assign targets_0_requests_5_valid = (gateways_4_ip && targets_0_ie_4);
  assign targets_0_requests_6_priority = gateways_5_priority;
  assign targets_0_requests_6_id = 5'h06;
  assign targets_0_requests_6_valid = (gateways_5_ip && targets_0_ie_5);
  assign targets_0_requests_7_priority = gateways_6_priority;
  assign targets_0_requests_7_id = 5'h07;
  assign targets_0_requests_7_valid = (gateways_6_ip && targets_0_ie_6);
  assign targets_0_requests_8_priority = gateways_7_priority;
  assign targets_0_requests_8_id = 5'h08;
  assign targets_0_requests_8_valid = (gateways_7_ip && targets_0_ie_7);
  assign targets_0_requests_9_priority = gateways_8_priority;
  assign targets_0_requests_9_id = 5'h09;
  assign targets_0_requests_9_valid = (gateways_8_ip && targets_0_ie_8);
  assign targets_0_requests_10_priority = gateways_9_priority;
  assign targets_0_requests_10_id = 5'h0a;
  assign targets_0_requests_10_valid = (gateways_9_ip && targets_0_ie_9);
  assign targets_0_requests_11_priority = gateways_10_priority;
  assign targets_0_requests_11_id = 5'h0b;
  assign targets_0_requests_11_valid = (gateways_10_ip && targets_0_ie_10);
  assign targets_0_requests_12_priority = gateways_11_priority;
  assign targets_0_requests_12_id = 5'h0c;
  assign targets_0_requests_12_valid = (gateways_11_ip && targets_0_ie_11);
  assign targets_0_requests_13_priority = gateways_12_priority;
  assign targets_0_requests_13_id = 5'h0d;
  assign targets_0_requests_13_valid = (gateways_12_ip && targets_0_ie_12);
  assign targets_0_requests_14_priority = gateways_13_priority;
  assign targets_0_requests_14_id = 5'h0e;
  assign targets_0_requests_14_valid = (gateways_13_ip && targets_0_ie_13);
  assign targets_0_requests_15_priority = gateways_14_priority;
  assign targets_0_requests_15_id = 5'h0f;
  assign targets_0_requests_15_valid = (gateways_14_ip && targets_0_ie_14);
  assign targets_0_requests_16_priority = gateways_15_priority;
  assign targets_0_requests_16_id = 5'h10;
  assign targets_0_requests_16_valid = (gateways_15_ip && targets_0_ie_15);
  assign targets_0_requests_17_priority = gateways_16_priority;
  assign targets_0_requests_17_id = 5'h11;
  assign targets_0_requests_17_valid = (gateways_16_ip && targets_0_ie_16);
  assign targets_0_requests_18_priority = gateways_17_priority;
  assign targets_0_requests_18_id = 5'h12;
  assign targets_0_requests_18_valid = (gateways_17_ip && targets_0_ie_17);
  assign targets_0_requests_19_priority = gateways_18_priority;
  assign targets_0_requests_19_id = 5'h13;
  assign targets_0_requests_19_valid = (gateways_18_ip && targets_0_ie_18);
  assign targets_0_requests_20_priority = gateways_19_priority;
  assign targets_0_requests_20_id = 5'h14;
  assign targets_0_requests_20_valid = (gateways_19_ip && targets_0_ie_19);
  assign targets_0_requests_21_priority = gateways_20_priority;
  assign targets_0_requests_21_id = 5'h15;
  assign targets_0_requests_21_valid = (gateways_20_ip && targets_0_ie_20);
  assign targets_0_requests_22_priority = gateways_21_priority;
  assign targets_0_requests_22_id = 5'h16;
  assign targets_0_requests_22_valid = (gateways_21_ip && targets_0_ie_21);
  assign targets_0_requests_23_priority = gateways_22_priority;
  assign targets_0_requests_23_id = 5'h17;
  assign targets_0_requests_23_valid = (gateways_22_ip && targets_0_ie_22);
  assign targets_0_requests_24_priority = gateways_23_priority;
  assign targets_0_requests_24_id = 5'h18;
  assign targets_0_requests_24_valid = (gateways_23_ip && targets_0_ie_23);
  assign targets_0_requests_25_priority = gateways_24_priority;
  assign targets_0_requests_25_id = 5'h19;
  assign targets_0_requests_25_valid = (gateways_24_ip && targets_0_ie_24);
  assign targets_0_requests_26_priority = gateways_25_priority;
  assign targets_0_requests_26_id = 5'h1a;
  assign targets_0_requests_26_valid = (gateways_25_ip && targets_0_ie_25);
  assign targets_0_requests_27_priority = gateways_26_priority;
  assign targets_0_requests_27_id = 5'h1b;
  assign targets_0_requests_27_valid = (gateways_26_ip && targets_0_ie_26);
  assign targets_0_requests_28_priority = gateways_27_priority;
  assign targets_0_requests_28_id = 5'h1c;
  assign targets_0_requests_28_valid = (gateways_27_ip && targets_0_ie_27);
  assign targets_0_requests_29_priority = gateways_28_priority;
  assign targets_0_requests_29_id = 5'h1d;
  assign targets_0_requests_29_valid = (gateways_28_ip && targets_0_ie_28);
  assign targets_0_requests_30_priority = gateways_29_priority;
  assign targets_0_requests_30_id = 5'h1e;
  assign targets_0_requests_30_valid = (gateways_29_ip && targets_0_ie_29);
  assign targets_0_requests_31_priority = gateways_30_priority;
  assign targets_0_requests_31_id = 5'h1f;
  assign targets_0_requests_31_valid = (gateways_30_ip && targets_0_ie_30);
  assign _zz_targets_0_bestRequest_id = ((! targets_0_requests_1_valid) || (targets_0_requests_0_valid && (targets_0_requests_1_priority <= targets_0_requests_0_priority)));
  assign _zz_targets_0_bestRequest_id_1 = (_zz_targets_0_bestRequest_id ? targets_0_requests_0_priority : targets_0_requests_1_priority);
  assign _zz_targets_0_bestRequest_id_2 = (_zz_targets_0_bestRequest_id ? targets_0_requests_0_valid : targets_0_requests_1_valid);
  assign _zz_targets_0_bestRequest_id_3 = ((! targets_0_requests_3_valid) || (targets_0_requests_2_valid && (targets_0_requests_3_priority <= targets_0_requests_2_priority)));
  assign _zz_targets_0_bestRequest_id_4 = (_zz_targets_0_bestRequest_id_3 ? targets_0_requests_2_priority : targets_0_requests_3_priority);
  assign _zz_targets_0_bestRequest_id_5 = (_zz_targets_0_bestRequest_id_3 ? targets_0_requests_2_valid : targets_0_requests_3_valid);
  assign _zz_targets_0_bestRequest_id_6 = ((! targets_0_requests_5_valid) || (targets_0_requests_4_valid && (targets_0_requests_5_priority <= targets_0_requests_4_priority)));
  assign _zz_targets_0_bestRequest_id_7 = (_zz_targets_0_bestRequest_id_6 ? targets_0_requests_4_priority : targets_0_requests_5_priority);
  assign _zz_targets_0_bestRequest_id_8 = (_zz_targets_0_bestRequest_id_6 ? targets_0_requests_4_valid : targets_0_requests_5_valid);
  assign _zz_targets_0_bestRequest_id_9 = ((! targets_0_requests_7_valid) || (targets_0_requests_6_valid && (targets_0_requests_7_priority <= targets_0_requests_6_priority)));
  assign _zz_targets_0_bestRequest_id_10 = (_zz_targets_0_bestRequest_id_9 ? targets_0_requests_6_priority : targets_0_requests_7_priority);
  assign _zz_targets_0_bestRequest_id_11 = (_zz_targets_0_bestRequest_id_9 ? targets_0_requests_6_valid : targets_0_requests_7_valid);
  assign _zz_targets_0_bestRequest_id_12 = ((! targets_0_requests_9_valid) || (targets_0_requests_8_valid && (targets_0_requests_9_priority <= targets_0_requests_8_priority)));
  assign _zz_targets_0_bestRequest_id_13 = (_zz_targets_0_bestRequest_id_12 ? targets_0_requests_8_priority : targets_0_requests_9_priority);
  assign _zz_targets_0_bestRequest_id_14 = (_zz_targets_0_bestRequest_id_12 ? targets_0_requests_8_valid : targets_0_requests_9_valid);
  assign _zz_targets_0_bestRequest_id_15 = ((! targets_0_requests_11_valid) || (targets_0_requests_10_valid && (targets_0_requests_11_priority <= targets_0_requests_10_priority)));
  assign _zz_targets_0_bestRequest_id_16 = (_zz_targets_0_bestRequest_id_15 ? targets_0_requests_10_priority : targets_0_requests_11_priority);
  assign _zz_targets_0_bestRequest_id_17 = (_zz_targets_0_bestRequest_id_15 ? targets_0_requests_10_valid : targets_0_requests_11_valid);
  assign _zz_targets_0_bestRequest_id_18 = ((! targets_0_requests_13_valid) || (targets_0_requests_12_valid && (targets_0_requests_13_priority <= targets_0_requests_12_priority)));
  assign _zz_targets_0_bestRequest_id_19 = (_zz_targets_0_bestRequest_id_18 ? targets_0_requests_12_priority : targets_0_requests_13_priority);
  assign _zz_targets_0_bestRequest_id_20 = (_zz_targets_0_bestRequest_id_18 ? targets_0_requests_12_valid : targets_0_requests_13_valid);
  assign _zz_targets_0_bestRequest_id_21 = ((! targets_0_requests_15_valid) || (targets_0_requests_14_valid && (targets_0_requests_15_priority <= targets_0_requests_14_priority)));
  assign _zz_targets_0_bestRequest_id_22 = (_zz_targets_0_bestRequest_id_21 ? targets_0_requests_14_priority : targets_0_requests_15_priority);
  assign _zz_targets_0_bestRequest_id_23 = (_zz_targets_0_bestRequest_id_21 ? targets_0_requests_14_valid : targets_0_requests_15_valid);
  assign _zz_targets_0_bestRequest_id_24 = ((! targets_0_requests_17_valid) || (targets_0_requests_16_valid && (targets_0_requests_17_priority <= targets_0_requests_16_priority)));
  assign _zz_targets_0_bestRequest_id_25 = (_zz_targets_0_bestRequest_id_24 ? targets_0_requests_16_priority : targets_0_requests_17_priority);
  assign _zz_targets_0_bestRequest_id_26 = (_zz_targets_0_bestRequest_id_24 ? targets_0_requests_16_valid : targets_0_requests_17_valid);
  assign _zz_targets_0_bestRequest_id_27 = ((! targets_0_requests_19_valid) || (targets_0_requests_18_valid && (targets_0_requests_19_priority <= targets_0_requests_18_priority)));
  assign _zz_targets_0_bestRequest_id_28 = (_zz_targets_0_bestRequest_id_27 ? targets_0_requests_18_priority : targets_0_requests_19_priority);
  assign _zz_targets_0_bestRequest_id_29 = (_zz_targets_0_bestRequest_id_27 ? targets_0_requests_18_valid : targets_0_requests_19_valid);
  assign _zz_targets_0_bestRequest_id_30 = ((! targets_0_requests_21_valid) || (targets_0_requests_20_valid && (targets_0_requests_21_priority <= targets_0_requests_20_priority)));
  assign _zz_targets_0_bestRequest_id_31 = (_zz_targets_0_bestRequest_id_30 ? targets_0_requests_20_priority : targets_0_requests_21_priority);
  assign _zz_targets_0_bestRequest_id_32 = (_zz_targets_0_bestRequest_id_30 ? targets_0_requests_20_valid : targets_0_requests_21_valid);
  assign _zz_targets_0_bestRequest_id_33 = ((! targets_0_requests_23_valid) || (targets_0_requests_22_valid && (targets_0_requests_23_priority <= targets_0_requests_22_priority)));
  assign _zz_targets_0_bestRequest_id_34 = (_zz_targets_0_bestRequest_id_33 ? targets_0_requests_22_priority : targets_0_requests_23_priority);
  assign _zz_targets_0_bestRequest_id_35 = (_zz_targets_0_bestRequest_id_33 ? targets_0_requests_22_valid : targets_0_requests_23_valid);
  assign _zz_targets_0_bestRequest_id_36 = ((! targets_0_requests_25_valid) || (targets_0_requests_24_valid && (targets_0_requests_25_priority <= targets_0_requests_24_priority)));
  assign _zz_targets_0_bestRequest_id_37 = (_zz_targets_0_bestRequest_id_36 ? targets_0_requests_24_priority : targets_0_requests_25_priority);
  assign _zz_targets_0_bestRequest_id_38 = (_zz_targets_0_bestRequest_id_36 ? targets_0_requests_24_valid : targets_0_requests_25_valid);
  assign _zz_targets_0_bestRequest_id_39 = ((! targets_0_requests_27_valid) || (targets_0_requests_26_valid && (targets_0_requests_27_priority <= targets_0_requests_26_priority)));
  assign _zz_targets_0_bestRequest_id_40 = (_zz_targets_0_bestRequest_id_39 ? targets_0_requests_26_priority : targets_0_requests_27_priority);
  assign _zz_targets_0_bestRequest_id_41 = (_zz_targets_0_bestRequest_id_39 ? targets_0_requests_26_valid : targets_0_requests_27_valid);
  assign _zz_targets_0_bestRequest_id_42 = ((! targets_0_requests_29_valid) || (targets_0_requests_28_valid && (targets_0_requests_29_priority <= targets_0_requests_28_priority)));
  assign _zz_targets_0_bestRequest_id_43 = (_zz_targets_0_bestRequest_id_42 ? targets_0_requests_28_priority : targets_0_requests_29_priority);
  assign _zz_targets_0_bestRequest_id_44 = (_zz_targets_0_bestRequest_id_42 ? targets_0_requests_28_valid : targets_0_requests_29_valid);
  assign _zz_targets_0_bestRequest_id_45 = ((! targets_0_requests_31_valid) || (targets_0_requests_30_valid && (targets_0_requests_31_priority <= targets_0_requests_30_priority)));
  assign _zz_targets_0_bestRequest_id_46 = (_zz_targets_0_bestRequest_id_45 ? targets_0_requests_30_priority : targets_0_requests_31_priority);
  assign _zz_targets_0_bestRequest_id_47 = (_zz_targets_0_bestRequest_id_45 ? targets_0_requests_30_valid : targets_0_requests_31_valid);
  assign _zz_targets_0_bestRequest_id_48 = ((! _zz_targets_0_bestRequest_id_5) || (_zz_targets_0_bestRequest_id_2 && (_zz_targets_0_bestRequest_id_4 <= _zz_targets_0_bestRequest_id_1)));
  assign _zz_targets_0_bestRequest_id_49 = (_zz_targets_0_bestRequest_id_48 ? _zz_targets_0_bestRequest_id_1 : _zz_targets_0_bestRequest_id_4);
  assign _zz_targets_0_bestRequest_id_50 = (_zz_targets_0_bestRequest_id_48 ? _zz_targets_0_bestRequest_id_2 : _zz_targets_0_bestRequest_id_5);
  assign _zz_targets_0_bestRequest_id_51 = ((! _zz_targets_0_bestRequest_id_11) || (_zz_targets_0_bestRequest_id_8 && (_zz_targets_0_bestRequest_id_10 <= _zz_targets_0_bestRequest_id_7)));
  assign _zz_targets_0_bestRequest_id_52 = (_zz_targets_0_bestRequest_id_51 ? _zz_targets_0_bestRequest_id_7 : _zz_targets_0_bestRequest_id_10);
  assign _zz_targets_0_bestRequest_id_53 = (_zz_targets_0_bestRequest_id_51 ? _zz_targets_0_bestRequest_id_8 : _zz_targets_0_bestRequest_id_11);
  assign _zz_targets_0_bestRequest_id_54 = ((! _zz_targets_0_bestRequest_id_17) || (_zz_targets_0_bestRequest_id_14 && (_zz_targets_0_bestRequest_id_16 <= _zz_targets_0_bestRequest_id_13)));
  assign _zz_targets_0_bestRequest_id_55 = (_zz_targets_0_bestRequest_id_54 ? _zz_targets_0_bestRequest_id_13 : _zz_targets_0_bestRequest_id_16);
  assign _zz_targets_0_bestRequest_id_56 = (_zz_targets_0_bestRequest_id_54 ? _zz_targets_0_bestRequest_id_14 : _zz_targets_0_bestRequest_id_17);
  assign _zz_targets_0_bestRequest_id_57 = ((! _zz_targets_0_bestRequest_id_23) || (_zz_targets_0_bestRequest_id_20 && (_zz_targets_0_bestRequest_id_22 <= _zz_targets_0_bestRequest_id_19)));
  assign _zz_targets_0_bestRequest_id_58 = (_zz_targets_0_bestRequest_id_57 ? _zz_targets_0_bestRequest_id_19 : _zz_targets_0_bestRequest_id_22);
  assign _zz_targets_0_bestRequest_id_59 = (_zz_targets_0_bestRequest_id_57 ? _zz_targets_0_bestRequest_id_20 : _zz_targets_0_bestRequest_id_23);
  assign _zz_targets_0_bestRequest_id_60 = ((! _zz_targets_0_bestRequest_id_29) || (_zz_targets_0_bestRequest_id_26 && (_zz_targets_0_bestRequest_id_28 <= _zz_targets_0_bestRequest_id_25)));
  assign _zz_targets_0_bestRequest_id_61 = (_zz_targets_0_bestRequest_id_60 ? _zz_targets_0_bestRequest_id_25 : _zz_targets_0_bestRequest_id_28);
  assign _zz_targets_0_bestRequest_id_62 = (_zz_targets_0_bestRequest_id_60 ? _zz_targets_0_bestRequest_id_26 : _zz_targets_0_bestRequest_id_29);
  assign _zz_targets_0_bestRequest_id_63 = ((! _zz_targets_0_bestRequest_id_35) || (_zz_targets_0_bestRequest_id_32 && (_zz_targets_0_bestRequest_id_34 <= _zz_targets_0_bestRequest_id_31)));
  assign _zz_targets_0_bestRequest_id_64 = (_zz_targets_0_bestRequest_id_63 ? _zz_targets_0_bestRequest_id_31 : _zz_targets_0_bestRequest_id_34);
  assign _zz_targets_0_bestRequest_id_65 = (_zz_targets_0_bestRequest_id_63 ? _zz_targets_0_bestRequest_id_32 : _zz_targets_0_bestRequest_id_35);
  assign _zz_targets_0_bestRequest_id_66 = ((! _zz_targets_0_bestRequest_id_41) || (_zz_targets_0_bestRequest_id_38 && (_zz_targets_0_bestRequest_id_40 <= _zz_targets_0_bestRequest_id_37)));
  assign _zz_targets_0_bestRequest_id_67 = (_zz_targets_0_bestRequest_id_66 ? _zz_targets_0_bestRequest_id_37 : _zz_targets_0_bestRequest_id_40);
  assign _zz_targets_0_bestRequest_id_68 = (_zz_targets_0_bestRequest_id_66 ? _zz_targets_0_bestRequest_id_38 : _zz_targets_0_bestRequest_id_41);
  assign _zz_targets_0_bestRequest_id_69 = ((! _zz_targets_0_bestRequest_id_47) || (_zz_targets_0_bestRequest_id_44 && (_zz_targets_0_bestRequest_id_46 <= _zz_targets_0_bestRequest_id_43)));
  assign _zz_targets_0_bestRequest_id_70 = (_zz_targets_0_bestRequest_id_69 ? _zz_targets_0_bestRequest_id_43 : _zz_targets_0_bestRequest_id_46);
  assign _zz_targets_0_bestRequest_id_71 = (_zz_targets_0_bestRequest_id_69 ? _zz_targets_0_bestRequest_id_44 : _zz_targets_0_bestRequest_id_47);
  assign _zz_targets_0_bestRequest_id_72 = ((! _zz_targets_0_bestRequest_id_53) || (_zz_targets_0_bestRequest_id_50 && (_zz_targets_0_bestRequest_id_52 <= _zz_targets_0_bestRequest_id_49)));
  assign _zz_targets_0_bestRequest_priority = (_zz_targets_0_bestRequest_id_72 ? _zz_targets_0_bestRequest_id_49 : _zz_targets_0_bestRequest_id_52);
  assign _zz_targets_0_bestRequest_id_73 = (_zz_targets_0_bestRequest_id_72 ? _zz_targets_0_bestRequest_id_50 : _zz_targets_0_bestRequest_id_53);
  assign _zz_targets_0_bestRequest_id_74 = ((! _zz_targets_0_bestRequest_id_59) || (_zz_targets_0_bestRequest_id_56 && (_zz_targets_0_bestRequest_id_58 <= _zz_targets_0_bestRequest_id_55)));
  assign _zz_targets_0_bestRequest_priority_1 = (_zz_targets_0_bestRequest_id_74 ? _zz_targets_0_bestRequest_id_55 : _zz_targets_0_bestRequest_id_58);
  assign _zz_targets_0_bestRequest_id_75 = (_zz_targets_0_bestRequest_id_74 ? _zz_targets_0_bestRequest_id_56 : _zz_targets_0_bestRequest_id_59);
  assign _zz_targets_0_bestRequest_id_76 = ((! _zz_targets_0_bestRequest_id_65) || (_zz_targets_0_bestRequest_id_62 && (_zz_targets_0_bestRequest_id_64 <= _zz_targets_0_bestRequest_id_61)));
  assign _zz_targets_0_bestRequest_priority_2 = (_zz_targets_0_bestRequest_id_76 ? _zz_targets_0_bestRequest_id_61 : _zz_targets_0_bestRequest_id_64);
  assign _zz_targets_0_bestRequest_id_77 = (_zz_targets_0_bestRequest_id_76 ? _zz_targets_0_bestRequest_id_62 : _zz_targets_0_bestRequest_id_65);
  assign _zz_targets_0_bestRequest_id_78 = ((! _zz_targets_0_bestRequest_id_71) || (_zz_targets_0_bestRequest_id_68 && (_zz_targets_0_bestRequest_id_70 <= _zz_targets_0_bestRequest_id_67)));
  assign _zz_targets_0_bestRequest_priority_3 = (_zz_targets_0_bestRequest_id_78 ? _zz_targets_0_bestRequest_id_67 : _zz_targets_0_bestRequest_id_70);
  assign _zz_targets_0_bestRequest_id_79 = (_zz_targets_0_bestRequest_id_78 ? _zz_targets_0_bestRequest_id_68 : _zz_targets_0_bestRequest_id_71);
  assign _zz_targets_0_bestRequest_id_80 = ((! _zz_targets_0_bestRequest_id_75) || (_zz_targets_0_bestRequest_id_73 && (_zz_targets_0_bestRequest_priority_1 <= _zz_targets_0_bestRequest_priority)));
  assign _zz_targets_0_bestRequest_priority_4 = (_zz_targets_0_bestRequest_id_80 ? _zz_targets_0_bestRequest_priority : _zz_targets_0_bestRequest_priority_1);
  assign _zz_targets_0_bestRequest_valid = (_zz_targets_0_bestRequest_id_80 ? _zz_targets_0_bestRequest_id_73 : _zz_targets_0_bestRequest_id_75);
  assign _zz_targets_0_bestRequest_id_81 = ((! _zz_targets_0_bestRequest_id_79) || (_zz_targets_0_bestRequest_id_77 && (_zz_targets_0_bestRequest_priority_3 <= _zz_targets_0_bestRequest_priority_2)));
  assign _zz_targets_0_bestRequest_priority_5 = (_zz_targets_0_bestRequest_id_81 ? _zz_targets_0_bestRequest_priority_2 : _zz_targets_0_bestRequest_priority_3);
  assign _zz_targets_0_bestRequest_valid_1 = (_zz_targets_0_bestRequest_id_81 ? _zz_targets_0_bestRequest_id_77 : _zz_targets_0_bestRequest_id_79);
  assign _zz_targets_0_bestRequest_priority_6 = ((! _zz_targets_0_bestRequest_valid_1) || (_zz_targets_0_bestRequest_valid && (_zz_targets_0_bestRequest_priority_5 <= _zz_targets_0_bestRequest_priority_4)));
  assign targets_0_iep = (targets_0_threshold < targets_0_bestRequest_priority);
  assign targets_0_claim = (targets_0_iep ? targets_0_bestRequest_id : 5'h00);
  assign targets_1_requests_0_priority = 2'b00;
  assign targets_1_requests_0_id = 5'h00;
  assign targets_1_requests_0_valid = 1'b1;
  assign targets_1_requests_1_priority = gateways_0_priority;
  assign targets_1_requests_1_id = 5'h01;
  assign targets_1_requests_1_valid = (gateways_0_ip && targets_1_ie_0);
  assign targets_1_requests_2_priority = gateways_1_priority;
  assign targets_1_requests_2_id = 5'h02;
  assign targets_1_requests_2_valid = (gateways_1_ip && targets_1_ie_1);
  assign targets_1_requests_3_priority = gateways_2_priority;
  assign targets_1_requests_3_id = 5'h03;
  assign targets_1_requests_3_valid = (gateways_2_ip && targets_1_ie_2);
  assign targets_1_requests_4_priority = gateways_3_priority;
  assign targets_1_requests_4_id = 5'h04;
  assign targets_1_requests_4_valid = (gateways_3_ip && targets_1_ie_3);
  assign targets_1_requests_5_priority = gateways_4_priority;
  assign targets_1_requests_5_id = 5'h05;
  assign targets_1_requests_5_valid = (gateways_4_ip && targets_1_ie_4);
  assign targets_1_requests_6_priority = gateways_5_priority;
  assign targets_1_requests_6_id = 5'h06;
  assign targets_1_requests_6_valid = (gateways_5_ip && targets_1_ie_5);
  assign targets_1_requests_7_priority = gateways_6_priority;
  assign targets_1_requests_7_id = 5'h07;
  assign targets_1_requests_7_valid = (gateways_6_ip && targets_1_ie_6);
  assign targets_1_requests_8_priority = gateways_7_priority;
  assign targets_1_requests_8_id = 5'h08;
  assign targets_1_requests_8_valid = (gateways_7_ip && targets_1_ie_7);
  assign targets_1_requests_9_priority = gateways_8_priority;
  assign targets_1_requests_9_id = 5'h09;
  assign targets_1_requests_9_valid = (gateways_8_ip && targets_1_ie_8);
  assign targets_1_requests_10_priority = gateways_9_priority;
  assign targets_1_requests_10_id = 5'h0a;
  assign targets_1_requests_10_valid = (gateways_9_ip && targets_1_ie_9);
  assign targets_1_requests_11_priority = gateways_10_priority;
  assign targets_1_requests_11_id = 5'h0b;
  assign targets_1_requests_11_valid = (gateways_10_ip && targets_1_ie_10);
  assign targets_1_requests_12_priority = gateways_11_priority;
  assign targets_1_requests_12_id = 5'h0c;
  assign targets_1_requests_12_valid = (gateways_11_ip && targets_1_ie_11);
  assign targets_1_requests_13_priority = gateways_12_priority;
  assign targets_1_requests_13_id = 5'h0d;
  assign targets_1_requests_13_valid = (gateways_12_ip && targets_1_ie_12);
  assign targets_1_requests_14_priority = gateways_13_priority;
  assign targets_1_requests_14_id = 5'h0e;
  assign targets_1_requests_14_valid = (gateways_13_ip && targets_1_ie_13);
  assign targets_1_requests_15_priority = gateways_14_priority;
  assign targets_1_requests_15_id = 5'h0f;
  assign targets_1_requests_15_valid = (gateways_14_ip && targets_1_ie_14);
  assign targets_1_requests_16_priority = gateways_15_priority;
  assign targets_1_requests_16_id = 5'h10;
  assign targets_1_requests_16_valid = (gateways_15_ip && targets_1_ie_15);
  assign targets_1_requests_17_priority = gateways_16_priority;
  assign targets_1_requests_17_id = 5'h11;
  assign targets_1_requests_17_valid = (gateways_16_ip && targets_1_ie_16);
  assign targets_1_requests_18_priority = gateways_17_priority;
  assign targets_1_requests_18_id = 5'h12;
  assign targets_1_requests_18_valid = (gateways_17_ip && targets_1_ie_17);
  assign targets_1_requests_19_priority = gateways_18_priority;
  assign targets_1_requests_19_id = 5'h13;
  assign targets_1_requests_19_valid = (gateways_18_ip && targets_1_ie_18);
  assign targets_1_requests_20_priority = gateways_19_priority;
  assign targets_1_requests_20_id = 5'h14;
  assign targets_1_requests_20_valid = (gateways_19_ip && targets_1_ie_19);
  assign targets_1_requests_21_priority = gateways_20_priority;
  assign targets_1_requests_21_id = 5'h15;
  assign targets_1_requests_21_valid = (gateways_20_ip && targets_1_ie_20);
  assign targets_1_requests_22_priority = gateways_21_priority;
  assign targets_1_requests_22_id = 5'h16;
  assign targets_1_requests_22_valid = (gateways_21_ip && targets_1_ie_21);
  assign targets_1_requests_23_priority = gateways_22_priority;
  assign targets_1_requests_23_id = 5'h17;
  assign targets_1_requests_23_valid = (gateways_22_ip && targets_1_ie_22);
  assign targets_1_requests_24_priority = gateways_23_priority;
  assign targets_1_requests_24_id = 5'h18;
  assign targets_1_requests_24_valid = (gateways_23_ip && targets_1_ie_23);
  assign targets_1_requests_25_priority = gateways_24_priority;
  assign targets_1_requests_25_id = 5'h19;
  assign targets_1_requests_25_valid = (gateways_24_ip && targets_1_ie_24);
  assign targets_1_requests_26_priority = gateways_25_priority;
  assign targets_1_requests_26_id = 5'h1a;
  assign targets_1_requests_26_valid = (gateways_25_ip && targets_1_ie_25);
  assign targets_1_requests_27_priority = gateways_26_priority;
  assign targets_1_requests_27_id = 5'h1b;
  assign targets_1_requests_27_valid = (gateways_26_ip && targets_1_ie_26);
  assign targets_1_requests_28_priority = gateways_27_priority;
  assign targets_1_requests_28_id = 5'h1c;
  assign targets_1_requests_28_valid = (gateways_27_ip && targets_1_ie_27);
  assign targets_1_requests_29_priority = gateways_28_priority;
  assign targets_1_requests_29_id = 5'h1d;
  assign targets_1_requests_29_valid = (gateways_28_ip && targets_1_ie_28);
  assign targets_1_requests_30_priority = gateways_29_priority;
  assign targets_1_requests_30_id = 5'h1e;
  assign targets_1_requests_30_valid = (gateways_29_ip && targets_1_ie_29);
  assign targets_1_requests_31_priority = gateways_30_priority;
  assign targets_1_requests_31_id = 5'h1f;
  assign targets_1_requests_31_valid = (gateways_30_ip && targets_1_ie_30);
  assign _zz_targets_1_bestRequest_id = ((! targets_1_requests_1_valid) || (targets_1_requests_0_valid && (targets_1_requests_1_priority <= targets_1_requests_0_priority)));
  assign _zz_targets_1_bestRequest_id_1 = (_zz_targets_1_bestRequest_id ? targets_1_requests_0_priority : targets_1_requests_1_priority);
  assign _zz_targets_1_bestRequest_id_2 = (_zz_targets_1_bestRequest_id ? targets_1_requests_0_valid : targets_1_requests_1_valid);
  assign _zz_targets_1_bestRequest_id_3 = ((! targets_1_requests_3_valid) || (targets_1_requests_2_valid && (targets_1_requests_3_priority <= targets_1_requests_2_priority)));
  assign _zz_targets_1_bestRequest_id_4 = (_zz_targets_1_bestRequest_id_3 ? targets_1_requests_2_priority : targets_1_requests_3_priority);
  assign _zz_targets_1_bestRequest_id_5 = (_zz_targets_1_bestRequest_id_3 ? targets_1_requests_2_valid : targets_1_requests_3_valid);
  assign _zz_targets_1_bestRequest_id_6 = ((! targets_1_requests_5_valid) || (targets_1_requests_4_valid && (targets_1_requests_5_priority <= targets_1_requests_4_priority)));
  assign _zz_targets_1_bestRequest_id_7 = (_zz_targets_1_bestRequest_id_6 ? targets_1_requests_4_priority : targets_1_requests_5_priority);
  assign _zz_targets_1_bestRequest_id_8 = (_zz_targets_1_bestRequest_id_6 ? targets_1_requests_4_valid : targets_1_requests_5_valid);
  assign _zz_targets_1_bestRequest_id_9 = ((! targets_1_requests_7_valid) || (targets_1_requests_6_valid && (targets_1_requests_7_priority <= targets_1_requests_6_priority)));
  assign _zz_targets_1_bestRequest_id_10 = (_zz_targets_1_bestRequest_id_9 ? targets_1_requests_6_priority : targets_1_requests_7_priority);
  assign _zz_targets_1_bestRequest_id_11 = (_zz_targets_1_bestRequest_id_9 ? targets_1_requests_6_valid : targets_1_requests_7_valid);
  assign _zz_targets_1_bestRequest_id_12 = ((! targets_1_requests_9_valid) || (targets_1_requests_8_valid && (targets_1_requests_9_priority <= targets_1_requests_8_priority)));
  assign _zz_targets_1_bestRequest_id_13 = (_zz_targets_1_bestRequest_id_12 ? targets_1_requests_8_priority : targets_1_requests_9_priority);
  assign _zz_targets_1_bestRequest_id_14 = (_zz_targets_1_bestRequest_id_12 ? targets_1_requests_8_valid : targets_1_requests_9_valid);
  assign _zz_targets_1_bestRequest_id_15 = ((! targets_1_requests_11_valid) || (targets_1_requests_10_valid && (targets_1_requests_11_priority <= targets_1_requests_10_priority)));
  assign _zz_targets_1_bestRequest_id_16 = (_zz_targets_1_bestRequest_id_15 ? targets_1_requests_10_priority : targets_1_requests_11_priority);
  assign _zz_targets_1_bestRequest_id_17 = (_zz_targets_1_bestRequest_id_15 ? targets_1_requests_10_valid : targets_1_requests_11_valid);
  assign _zz_targets_1_bestRequest_id_18 = ((! targets_1_requests_13_valid) || (targets_1_requests_12_valid && (targets_1_requests_13_priority <= targets_1_requests_12_priority)));
  assign _zz_targets_1_bestRequest_id_19 = (_zz_targets_1_bestRequest_id_18 ? targets_1_requests_12_priority : targets_1_requests_13_priority);
  assign _zz_targets_1_bestRequest_id_20 = (_zz_targets_1_bestRequest_id_18 ? targets_1_requests_12_valid : targets_1_requests_13_valid);
  assign _zz_targets_1_bestRequest_id_21 = ((! targets_1_requests_15_valid) || (targets_1_requests_14_valid && (targets_1_requests_15_priority <= targets_1_requests_14_priority)));
  assign _zz_targets_1_bestRequest_id_22 = (_zz_targets_1_bestRequest_id_21 ? targets_1_requests_14_priority : targets_1_requests_15_priority);
  assign _zz_targets_1_bestRequest_id_23 = (_zz_targets_1_bestRequest_id_21 ? targets_1_requests_14_valid : targets_1_requests_15_valid);
  assign _zz_targets_1_bestRequest_id_24 = ((! targets_1_requests_17_valid) || (targets_1_requests_16_valid && (targets_1_requests_17_priority <= targets_1_requests_16_priority)));
  assign _zz_targets_1_bestRequest_id_25 = (_zz_targets_1_bestRequest_id_24 ? targets_1_requests_16_priority : targets_1_requests_17_priority);
  assign _zz_targets_1_bestRequest_id_26 = (_zz_targets_1_bestRequest_id_24 ? targets_1_requests_16_valid : targets_1_requests_17_valid);
  assign _zz_targets_1_bestRequest_id_27 = ((! targets_1_requests_19_valid) || (targets_1_requests_18_valid && (targets_1_requests_19_priority <= targets_1_requests_18_priority)));
  assign _zz_targets_1_bestRequest_id_28 = (_zz_targets_1_bestRequest_id_27 ? targets_1_requests_18_priority : targets_1_requests_19_priority);
  assign _zz_targets_1_bestRequest_id_29 = (_zz_targets_1_bestRequest_id_27 ? targets_1_requests_18_valid : targets_1_requests_19_valid);
  assign _zz_targets_1_bestRequest_id_30 = ((! targets_1_requests_21_valid) || (targets_1_requests_20_valid && (targets_1_requests_21_priority <= targets_1_requests_20_priority)));
  assign _zz_targets_1_bestRequest_id_31 = (_zz_targets_1_bestRequest_id_30 ? targets_1_requests_20_priority : targets_1_requests_21_priority);
  assign _zz_targets_1_bestRequest_id_32 = (_zz_targets_1_bestRequest_id_30 ? targets_1_requests_20_valid : targets_1_requests_21_valid);
  assign _zz_targets_1_bestRequest_id_33 = ((! targets_1_requests_23_valid) || (targets_1_requests_22_valid && (targets_1_requests_23_priority <= targets_1_requests_22_priority)));
  assign _zz_targets_1_bestRequest_id_34 = (_zz_targets_1_bestRequest_id_33 ? targets_1_requests_22_priority : targets_1_requests_23_priority);
  assign _zz_targets_1_bestRequest_id_35 = (_zz_targets_1_bestRequest_id_33 ? targets_1_requests_22_valid : targets_1_requests_23_valid);
  assign _zz_targets_1_bestRequest_id_36 = ((! targets_1_requests_25_valid) || (targets_1_requests_24_valid && (targets_1_requests_25_priority <= targets_1_requests_24_priority)));
  assign _zz_targets_1_bestRequest_id_37 = (_zz_targets_1_bestRequest_id_36 ? targets_1_requests_24_priority : targets_1_requests_25_priority);
  assign _zz_targets_1_bestRequest_id_38 = (_zz_targets_1_bestRequest_id_36 ? targets_1_requests_24_valid : targets_1_requests_25_valid);
  assign _zz_targets_1_bestRequest_id_39 = ((! targets_1_requests_27_valid) || (targets_1_requests_26_valid && (targets_1_requests_27_priority <= targets_1_requests_26_priority)));
  assign _zz_targets_1_bestRequest_id_40 = (_zz_targets_1_bestRequest_id_39 ? targets_1_requests_26_priority : targets_1_requests_27_priority);
  assign _zz_targets_1_bestRequest_id_41 = (_zz_targets_1_bestRequest_id_39 ? targets_1_requests_26_valid : targets_1_requests_27_valid);
  assign _zz_targets_1_bestRequest_id_42 = ((! targets_1_requests_29_valid) || (targets_1_requests_28_valid && (targets_1_requests_29_priority <= targets_1_requests_28_priority)));
  assign _zz_targets_1_bestRequest_id_43 = (_zz_targets_1_bestRequest_id_42 ? targets_1_requests_28_priority : targets_1_requests_29_priority);
  assign _zz_targets_1_bestRequest_id_44 = (_zz_targets_1_bestRequest_id_42 ? targets_1_requests_28_valid : targets_1_requests_29_valid);
  assign _zz_targets_1_bestRequest_id_45 = ((! targets_1_requests_31_valid) || (targets_1_requests_30_valid && (targets_1_requests_31_priority <= targets_1_requests_30_priority)));
  assign _zz_targets_1_bestRequest_id_46 = (_zz_targets_1_bestRequest_id_45 ? targets_1_requests_30_priority : targets_1_requests_31_priority);
  assign _zz_targets_1_bestRequest_id_47 = (_zz_targets_1_bestRequest_id_45 ? targets_1_requests_30_valid : targets_1_requests_31_valid);
  assign _zz_targets_1_bestRequest_id_48 = ((! _zz_targets_1_bestRequest_id_5) || (_zz_targets_1_bestRequest_id_2 && (_zz_targets_1_bestRequest_id_4 <= _zz_targets_1_bestRequest_id_1)));
  assign _zz_targets_1_bestRequest_id_49 = (_zz_targets_1_bestRequest_id_48 ? _zz_targets_1_bestRequest_id_1 : _zz_targets_1_bestRequest_id_4);
  assign _zz_targets_1_bestRequest_id_50 = (_zz_targets_1_bestRequest_id_48 ? _zz_targets_1_bestRequest_id_2 : _zz_targets_1_bestRequest_id_5);
  assign _zz_targets_1_bestRequest_id_51 = ((! _zz_targets_1_bestRequest_id_11) || (_zz_targets_1_bestRequest_id_8 && (_zz_targets_1_bestRequest_id_10 <= _zz_targets_1_bestRequest_id_7)));
  assign _zz_targets_1_bestRequest_id_52 = (_zz_targets_1_bestRequest_id_51 ? _zz_targets_1_bestRequest_id_7 : _zz_targets_1_bestRequest_id_10);
  assign _zz_targets_1_bestRequest_id_53 = (_zz_targets_1_bestRequest_id_51 ? _zz_targets_1_bestRequest_id_8 : _zz_targets_1_bestRequest_id_11);
  assign _zz_targets_1_bestRequest_id_54 = ((! _zz_targets_1_bestRequest_id_17) || (_zz_targets_1_bestRequest_id_14 && (_zz_targets_1_bestRequest_id_16 <= _zz_targets_1_bestRequest_id_13)));
  assign _zz_targets_1_bestRequest_id_55 = (_zz_targets_1_bestRequest_id_54 ? _zz_targets_1_bestRequest_id_13 : _zz_targets_1_bestRequest_id_16);
  assign _zz_targets_1_bestRequest_id_56 = (_zz_targets_1_bestRequest_id_54 ? _zz_targets_1_bestRequest_id_14 : _zz_targets_1_bestRequest_id_17);
  assign _zz_targets_1_bestRequest_id_57 = ((! _zz_targets_1_bestRequest_id_23) || (_zz_targets_1_bestRequest_id_20 && (_zz_targets_1_bestRequest_id_22 <= _zz_targets_1_bestRequest_id_19)));
  assign _zz_targets_1_bestRequest_id_58 = (_zz_targets_1_bestRequest_id_57 ? _zz_targets_1_bestRequest_id_19 : _zz_targets_1_bestRequest_id_22);
  assign _zz_targets_1_bestRequest_id_59 = (_zz_targets_1_bestRequest_id_57 ? _zz_targets_1_bestRequest_id_20 : _zz_targets_1_bestRequest_id_23);
  assign _zz_targets_1_bestRequest_id_60 = ((! _zz_targets_1_bestRequest_id_29) || (_zz_targets_1_bestRequest_id_26 && (_zz_targets_1_bestRequest_id_28 <= _zz_targets_1_bestRequest_id_25)));
  assign _zz_targets_1_bestRequest_id_61 = (_zz_targets_1_bestRequest_id_60 ? _zz_targets_1_bestRequest_id_25 : _zz_targets_1_bestRequest_id_28);
  assign _zz_targets_1_bestRequest_id_62 = (_zz_targets_1_bestRequest_id_60 ? _zz_targets_1_bestRequest_id_26 : _zz_targets_1_bestRequest_id_29);
  assign _zz_targets_1_bestRequest_id_63 = ((! _zz_targets_1_bestRequest_id_35) || (_zz_targets_1_bestRequest_id_32 && (_zz_targets_1_bestRequest_id_34 <= _zz_targets_1_bestRequest_id_31)));
  assign _zz_targets_1_bestRequest_id_64 = (_zz_targets_1_bestRequest_id_63 ? _zz_targets_1_bestRequest_id_31 : _zz_targets_1_bestRequest_id_34);
  assign _zz_targets_1_bestRequest_id_65 = (_zz_targets_1_bestRequest_id_63 ? _zz_targets_1_bestRequest_id_32 : _zz_targets_1_bestRequest_id_35);
  assign _zz_targets_1_bestRequest_id_66 = ((! _zz_targets_1_bestRequest_id_41) || (_zz_targets_1_bestRequest_id_38 && (_zz_targets_1_bestRequest_id_40 <= _zz_targets_1_bestRequest_id_37)));
  assign _zz_targets_1_bestRequest_id_67 = (_zz_targets_1_bestRequest_id_66 ? _zz_targets_1_bestRequest_id_37 : _zz_targets_1_bestRequest_id_40);
  assign _zz_targets_1_bestRequest_id_68 = (_zz_targets_1_bestRequest_id_66 ? _zz_targets_1_bestRequest_id_38 : _zz_targets_1_bestRequest_id_41);
  assign _zz_targets_1_bestRequest_id_69 = ((! _zz_targets_1_bestRequest_id_47) || (_zz_targets_1_bestRequest_id_44 && (_zz_targets_1_bestRequest_id_46 <= _zz_targets_1_bestRequest_id_43)));
  assign _zz_targets_1_bestRequest_id_70 = (_zz_targets_1_bestRequest_id_69 ? _zz_targets_1_bestRequest_id_43 : _zz_targets_1_bestRequest_id_46);
  assign _zz_targets_1_bestRequest_id_71 = (_zz_targets_1_bestRequest_id_69 ? _zz_targets_1_bestRequest_id_44 : _zz_targets_1_bestRequest_id_47);
  assign _zz_targets_1_bestRequest_id_72 = ((! _zz_targets_1_bestRequest_id_53) || (_zz_targets_1_bestRequest_id_50 && (_zz_targets_1_bestRequest_id_52 <= _zz_targets_1_bestRequest_id_49)));
  assign _zz_targets_1_bestRequest_priority = (_zz_targets_1_bestRequest_id_72 ? _zz_targets_1_bestRequest_id_49 : _zz_targets_1_bestRequest_id_52);
  assign _zz_targets_1_bestRequest_id_73 = (_zz_targets_1_bestRequest_id_72 ? _zz_targets_1_bestRequest_id_50 : _zz_targets_1_bestRequest_id_53);
  assign _zz_targets_1_bestRequest_id_74 = ((! _zz_targets_1_bestRequest_id_59) || (_zz_targets_1_bestRequest_id_56 && (_zz_targets_1_bestRequest_id_58 <= _zz_targets_1_bestRequest_id_55)));
  assign _zz_targets_1_bestRequest_priority_1 = (_zz_targets_1_bestRequest_id_74 ? _zz_targets_1_bestRequest_id_55 : _zz_targets_1_bestRequest_id_58);
  assign _zz_targets_1_bestRequest_id_75 = (_zz_targets_1_bestRequest_id_74 ? _zz_targets_1_bestRequest_id_56 : _zz_targets_1_bestRequest_id_59);
  assign _zz_targets_1_bestRequest_id_76 = ((! _zz_targets_1_bestRequest_id_65) || (_zz_targets_1_bestRequest_id_62 && (_zz_targets_1_bestRequest_id_64 <= _zz_targets_1_bestRequest_id_61)));
  assign _zz_targets_1_bestRequest_priority_2 = (_zz_targets_1_bestRequest_id_76 ? _zz_targets_1_bestRequest_id_61 : _zz_targets_1_bestRequest_id_64);
  assign _zz_targets_1_bestRequest_id_77 = (_zz_targets_1_bestRequest_id_76 ? _zz_targets_1_bestRequest_id_62 : _zz_targets_1_bestRequest_id_65);
  assign _zz_targets_1_bestRequest_id_78 = ((! _zz_targets_1_bestRequest_id_71) || (_zz_targets_1_bestRequest_id_68 && (_zz_targets_1_bestRequest_id_70 <= _zz_targets_1_bestRequest_id_67)));
  assign _zz_targets_1_bestRequest_priority_3 = (_zz_targets_1_bestRequest_id_78 ? _zz_targets_1_bestRequest_id_67 : _zz_targets_1_bestRequest_id_70);
  assign _zz_targets_1_bestRequest_id_79 = (_zz_targets_1_bestRequest_id_78 ? _zz_targets_1_bestRequest_id_68 : _zz_targets_1_bestRequest_id_71);
  assign _zz_targets_1_bestRequest_id_80 = ((! _zz_targets_1_bestRequest_id_75) || (_zz_targets_1_bestRequest_id_73 && (_zz_targets_1_bestRequest_priority_1 <= _zz_targets_1_bestRequest_priority)));
  assign _zz_targets_1_bestRequest_priority_4 = (_zz_targets_1_bestRequest_id_80 ? _zz_targets_1_bestRequest_priority : _zz_targets_1_bestRequest_priority_1);
  assign _zz_targets_1_bestRequest_valid = (_zz_targets_1_bestRequest_id_80 ? _zz_targets_1_bestRequest_id_73 : _zz_targets_1_bestRequest_id_75);
  assign _zz_targets_1_bestRequest_id_81 = ((! _zz_targets_1_bestRequest_id_79) || (_zz_targets_1_bestRequest_id_77 && (_zz_targets_1_bestRequest_priority_3 <= _zz_targets_1_bestRequest_priority_2)));
  assign _zz_targets_1_bestRequest_priority_5 = (_zz_targets_1_bestRequest_id_81 ? _zz_targets_1_bestRequest_priority_2 : _zz_targets_1_bestRequest_priority_3);
  assign _zz_targets_1_bestRequest_valid_1 = (_zz_targets_1_bestRequest_id_81 ? _zz_targets_1_bestRequest_id_77 : _zz_targets_1_bestRequest_id_79);
  assign _zz_targets_1_bestRequest_priority_6 = ((! _zz_targets_1_bestRequest_valid_1) || (_zz_targets_1_bestRequest_valid && (_zz_targets_1_bestRequest_priority_5 <= _zz_targets_1_bestRequest_priority_4)));
  assign targets_1_iep = (targets_1_threshold < targets_1_bestRequest_priority);
  assign targets_1_claim = (targets_1_iep ? targets_1_bestRequest_id : 5'h00);
  assign io_targets = {targets_1_iep,targets_0_iep};
  assign bus_readErrorFlag = 1'b0;
  assign bus_writeErrorFlag = 1'b0;
  always @(*) begin
    bus_readHaltRequest = 1'b0;
    if(when_PlicMapper_l122) begin
      bus_readHaltRequest = 1'b1;
    end
  end

  assign bus_writeHaltRequest = 1'b0;
  assign bus_writeOccur = (bus_writeJoinEvent_valid && bus_writeJoinEvent_ready);
  assign bus_writeJoinEvent_valid = (io_bus_aw_valid && io_bus_w_valid);
  assign io_bus_aw_ready = bus_writeOccur;
  assign io_bus_w_ready = bus_writeOccur;
  assign bus_writeJoinEvent_translated_valid = bus_writeJoinEvent_valid;
  assign bus_writeJoinEvent_ready = bus_writeJoinEvent_translated_ready;
  assign bus_writeJoinEvent_translated_payload_resp = bus_writeRsp_resp;
  assign _zz_bus_writeJoinEvent_translated_ready = (! bus_writeHaltRequest);
  assign bus_writeJoinEvent_translated_ready = (_zz_bus_writeJoinEvent_translated_ready_1 && _zz_bus_writeJoinEvent_translated_ready);
  assign _zz_bus_writeJoinEvent_translated_ready_1 = (! _zz_io_bus_b_valid_1);
  assign _zz_io_bus_b_valid = _zz_io_bus_b_valid_1;
  assign io_bus_b_valid = _zz_io_bus_b_valid;
  assign io_bus_b_payload_resp = _zz_io_bus_b_payload_resp;
  assign bus_readDataStage_fire = (bus_readDataStage_valid && bus_readDataStage_ready);
  assign io_bus_ar_ready = (! io_bus_ar_rValid);
  assign bus_readDataStage_valid = io_bus_ar_rValid;
  assign bus_readDataStage_payload_addr = io_bus_ar_rData_addr;
  assign bus_readDataStage_payload_prot = io_bus_ar_rData_prot;
  assign _zz_io_bus_r_valid = (! bus_readHaltRequest);
  assign bus_readDataStage_ready = (io_bus_r_ready && _zz_io_bus_r_valid);
  assign io_bus_r_valid = (bus_readDataStage_valid && _zz_io_bus_r_valid);
  assign io_bus_r_payload_data = bus_readRsp_data;
  assign io_bus_r_payload_resp = bus_readRsp_resp;
  always @(*) begin
    if(bus_writeErrorFlag) begin
      bus_writeRsp_resp = 2'b10;
    end else begin
      bus_writeRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    if(bus_readErrorFlag) begin
      bus_readRsp_resp = 2'b10;
    end else begin
      bus_readRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    bus_readRsp_data = 32'h00000000;
    case(bus_readAddressMasked)
      22'h000004 : begin
        bus_readRsp_data[1 : 0] = gateways_0_priority;
      end
      22'h001000 : begin
        bus_readRsp_data[1 : 1] = gateways_0_ip;
        bus_readRsp_data[2 : 2] = gateways_1_ip;
        bus_readRsp_data[3 : 3] = gateways_2_ip;
        bus_readRsp_data[4 : 4] = gateways_3_ip;
        bus_readRsp_data[5 : 5] = gateways_4_ip;
        bus_readRsp_data[6 : 6] = gateways_5_ip;
        bus_readRsp_data[7 : 7] = gateways_6_ip;
        bus_readRsp_data[8 : 8] = gateways_7_ip;
        bus_readRsp_data[9 : 9] = gateways_8_ip;
        bus_readRsp_data[10 : 10] = gateways_9_ip;
        bus_readRsp_data[11 : 11] = gateways_10_ip;
        bus_readRsp_data[12 : 12] = gateways_11_ip;
        bus_readRsp_data[13 : 13] = gateways_12_ip;
        bus_readRsp_data[14 : 14] = gateways_13_ip;
        bus_readRsp_data[15 : 15] = gateways_14_ip;
        bus_readRsp_data[16 : 16] = gateways_15_ip;
        bus_readRsp_data[17 : 17] = gateways_16_ip;
        bus_readRsp_data[18 : 18] = gateways_17_ip;
        bus_readRsp_data[19 : 19] = gateways_18_ip;
        bus_readRsp_data[20 : 20] = gateways_19_ip;
        bus_readRsp_data[21 : 21] = gateways_20_ip;
        bus_readRsp_data[22 : 22] = gateways_21_ip;
        bus_readRsp_data[23 : 23] = gateways_22_ip;
        bus_readRsp_data[24 : 24] = gateways_23_ip;
        bus_readRsp_data[25 : 25] = gateways_24_ip;
        bus_readRsp_data[26 : 26] = gateways_25_ip;
        bus_readRsp_data[27 : 27] = gateways_26_ip;
        bus_readRsp_data[28 : 28] = gateways_27_ip;
        bus_readRsp_data[29 : 29] = gateways_28_ip;
        bus_readRsp_data[30 : 30] = gateways_29_ip;
        bus_readRsp_data[31 : 31] = gateways_30_ip;
      end
      22'h000008 : begin
        bus_readRsp_data[1 : 0] = gateways_1_priority;
      end
      22'h00000c : begin
        bus_readRsp_data[1 : 0] = gateways_2_priority;
      end
      22'h000010 : begin
        bus_readRsp_data[1 : 0] = gateways_3_priority;
      end
      22'h000014 : begin
        bus_readRsp_data[1 : 0] = gateways_4_priority;
      end
      22'h000018 : begin
        bus_readRsp_data[1 : 0] = gateways_5_priority;
      end
      22'h00001c : begin
        bus_readRsp_data[1 : 0] = gateways_6_priority;
      end
      22'h000020 : begin
        bus_readRsp_data[1 : 0] = gateways_7_priority;
      end
      22'h000024 : begin
        bus_readRsp_data[1 : 0] = gateways_8_priority;
      end
      22'h000028 : begin
        bus_readRsp_data[1 : 0] = gateways_9_priority;
      end
      22'h00002c : begin
        bus_readRsp_data[1 : 0] = gateways_10_priority;
      end
      22'h000030 : begin
        bus_readRsp_data[1 : 0] = gateways_11_priority;
      end
      22'h000034 : begin
        bus_readRsp_data[1 : 0] = gateways_12_priority;
      end
      22'h000038 : begin
        bus_readRsp_data[1 : 0] = gateways_13_priority;
      end
      22'h00003c : begin
        bus_readRsp_data[1 : 0] = gateways_14_priority;
      end
      22'h000040 : begin
        bus_readRsp_data[1 : 0] = gateways_15_priority;
      end
      22'h000044 : begin
        bus_readRsp_data[1 : 0] = gateways_16_priority;
      end
      22'h000048 : begin
        bus_readRsp_data[1 : 0] = gateways_17_priority;
      end
      22'h00004c : begin
        bus_readRsp_data[1 : 0] = gateways_18_priority;
      end
      22'h000050 : begin
        bus_readRsp_data[1 : 0] = gateways_19_priority;
      end
      22'h000054 : begin
        bus_readRsp_data[1 : 0] = gateways_20_priority;
      end
      22'h000058 : begin
        bus_readRsp_data[1 : 0] = gateways_21_priority;
      end
      22'h00005c : begin
        bus_readRsp_data[1 : 0] = gateways_22_priority;
      end
      22'h000060 : begin
        bus_readRsp_data[1 : 0] = gateways_23_priority;
      end
      22'h000064 : begin
        bus_readRsp_data[1 : 0] = gateways_24_priority;
      end
      22'h000068 : begin
        bus_readRsp_data[1 : 0] = gateways_25_priority;
      end
      22'h00006c : begin
        bus_readRsp_data[1 : 0] = gateways_26_priority;
      end
      22'h000070 : begin
        bus_readRsp_data[1 : 0] = gateways_27_priority;
      end
      22'h000074 : begin
        bus_readRsp_data[1 : 0] = gateways_28_priority;
      end
      22'h000078 : begin
        bus_readRsp_data[1 : 0] = gateways_29_priority;
      end
      22'h00007c : begin
        bus_readRsp_data[1 : 0] = gateways_30_priority;
      end
      22'h200000 : begin
        bus_readRsp_data[1 : 0] = targets_0_threshold;
      end
      22'h200004 : begin
        bus_readRsp_data[4 : 0] = targets_0_claim;
      end
      22'h002000 : begin
        bus_readRsp_data[1 : 1] = targets_0_ie_0;
        bus_readRsp_data[2 : 2] = targets_0_ie_1;
        bus_readRsp_data[3 : 3] = targets_0_ie_2;
        bus_readRsp_data[4 : 4] = targets_0_ie_3;
        bus_readRsp_data[5 : 5] = targets_0_ie_4;
        bus_readRsp_data[6 : 6] = targets_0_ie_5;
        bus_readRsp_data[7 : 7] = targets_0_ie_6;
        bus_readRsp_data[8 : 8] = targets_0_ie_7;
        bus_readRsp_data[9 : 9] = targets_0_ie_8;
        bus_readRsp_data[10 : 10] = targets_0_ie_9;
        bus_readRsp_data[11 : 11] = targets_0_ie_10;
        bus_readRsp_data[12 : 12] = targets_0_ie_11;
        bus_readRsp_data[13 : 13] = targets_0_ie_12;
        bus_readRsp_data[14 : 14] = targets_0_ie_13;
        bus_readRsp_data[15 : 15] = targets_0_ie_14;
        bus_readRsp_data[16 : 16] = targets_0_ie_15;
        bus_readRsp_data[17 : 17] = targets_0_ie_16;
        bus_readRsp_data[18 : 18] = targets_0_ie_17;
        bus_readRsp_data[19 : 19] = targets_0_ie_18;
        bus_readRsp_data[20 : 20] = targets_0_ie_19;
        bus_readRsp_data[21 : 21] = targets_0_ie_20;
        bus_readRsp_data[22 : 22] = targets_0_ie_21;
        bus_readRsp_data[23 : 23] = targets_0_ie_22;
        bus_readRsp_data[24 : 24] = targets_0_ie_23;
        bus_readRsp_data[25 : 25] = targets_0_ie_24;
        bus_readRsp_data[26 : 26] = targets_0_ie_25;
        bus_readRsp_data[27 : 27] = targets_0_ie_26;
        bus_readRsp_data[28 : 28] = targets_0_ie_27;
        bus_readRsp_data[29 : 29] = targets_0_ie_28;
        bus_readRsp_data[30 : 30] = targets_0_ie_29;
        bus_readRsp_data[31 : 31] = targets_0_ie_30;
      end
      22'h201000 : begin
        bus_readRsp_data[1 : 0] = targets_1_threshold;
      end
      22'h201004 : begin
        bus_readRsp_data[4 : 0] = targets_1_claim;
      end
      22'h002080 : begin
        bus_readRsp_data[1 : 1] = targets_1_ie_0;
        bus_readRsp_data[2 : 2] = targets_1_ie_1;
        bus_readRsp_data[3 : 3] = targets_1_ie_2;
        bus_readRsp_data[4 : 4] = targets_1_ie_3;
        bus_readRsp_data[5 : 5] = targets_1_ie_4;
        bus_readRsp_data[6 : 6] = targets_1_ie_5;
        bus_readRsp_data[7 : 7] = targets_1_ie_6;
        bus_readRsp_data[8 : 8] = targets_1_ie_7;
        bus_readRsp_data[9 : 9] = targets_1_ie_8;
        bus_readRsp_data[10 : 10] = targets_1_ie_9;
        bus_readRsp_data[11 : 11] = targets_1_ie_10;
        bus_readRsp_data[12 : 12] = targets_1_ie_11;
        bus_readRsp_data[13 : 13] = targets_1_ie_12;
        bus_readRsp_data[14 : 14] = targets_1_ie_13;
        bus_readRsp_data[15 : 15] = targets_1_ie_14;
        bus_readRsp_data[16 : 16] = targets_1_ie_15;
        bus_readRsp_data[17 : 17] = targets_1_ie_16;
        bus_readRsp_data[18 : 18] = targets_1_ie_17;
        bus_readRsp_data[19 : 19] = targets_1_ie_18;
        bus_readRsp_data[20 : 20] = targets_1_ie_19;
        bus_readRsp_data[21 : 21] = targets_1_ie_20;
        bus_readRsp_data[22 : 22] = targets_1_ie_21;
        bus_readRsp_data[23 : 23] = targets_1_ie_22;
        bus_readRsp_data[24 : 24] = targets_1_ie_23;
        bus_readRsp_data[25 : 25] = targets_1_ie_24;
        bus_readRsp_data[26 : 26] = targets_1_ie_25;
        bus_readRsp_data[27 : 27] = targets_1_ie_26;
        bus_readRsp_data[28 : 28] = targets_1_ie_27;
        bus_readRsp_data[29 : 29] = targets_1_ie_28;
        bus_readRsp_data[30 : 30] = targets_1_ie_29;
        bus_readRsp_data[31 : 31] = targets_1_ie_30;
      end
      default : begin
      end
    endcase
  end

  assign bus_readAddressMasked = (bus_readDataStage_payload_addr & (~ 22'h000003));
  assign bus_writeAddressMasked = (io_bus_aw_payload_addr & (~ 22'h000003));
  assign bus_readOccur = (io_bus_r_valid && io_bus_r_ready);
  assign gateways_0_priority = _zz_gateways_0_priority;
  assign gateways_1_priority = _zz_gateways_1_priority;
  assign gateways_2_priority = _zz_gateways_2_priority;
  assign gateways_3_priority = _zz_gateways_3_priority;
  assign gateways_4_priority = _zz_gateways_4_priority;
  assign gateways_5_priority = _zz_gateways_5_priority;
  assign gateways_6_priority = _zz_gateways_6_priority;
  assign gateways_7_priority = _zz_gateways_7_priority;
  assign gateways_8_priority = _zz_gateways_8_priority;
  assign gateways_9_priority = _zz_gateways_9_priority;
  assign gateways_10_priority = _zz_gateways_10_priority;
  assign gateways_11_priority = _zz_gateways_11_priority;
  assign gateways_12_priority = _zz_gateways_12_priority;
  assign gateways_13_priority = _zz_gateways_13_priority;
  assign gateways_14_priority = _zz_gateways_14_priority;
  assign gateways_15_priority = _zz_gateways_15_priority;
  assign gateways_16_priority = _zz_gateways_16_priority;
  assign gateways_17_priority = _zz_gateways_17_priority;
  assign gateways_18_priority = _zz_gateways_18_priority;
  assign gateways_19_priority = _zz_gateways_19_priority;
  assign gateways_20_priority = _zz_gateways_20_priority;
  assign gateways_21_priority = _zz_gateways_21_priority;
  assign gateways_22_priority = _zz_gateways_22_priority;
  assign gateways_23_priority = _zz_gateways_23_priority;
  assign gateways_24_priority = _zz_gateways_24_priority;
  assign gateways_25_priority = _zz_gateways_25_priority;
  assign gateways_26_priority = _zz_gateways_26_priority;
  assign gateways_27_priority = _zz_gateways_27_priority;
  assign gateways_28_priority = _zz_gateways_28_priority;
  assign gateways_29_priority = _zz_gateways_29_priority;
  assign gateways_30_priority = _zz_gateways_30_priority;
  always @(*) begin
    mapping_claim_valid = 1'b0;
    case(bus_readAddressMasked)
      22'h200004 : begin
        if(bus_readOccur) begin
          mapping_claim_valid = 1'b1;
        end
      end
      22'h201004 : begin
        if(bus_readOccur) begin
          mapping_claim_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mapping_claim_payload = 5'bxxxxx;
    case(bus_readAddressMasked)
      22'h200004 : begin
        if(bus_readOccur) begin
          mapping_claim_payload = targets_0_claim;
        end
      end
      22'h201004 : begin
        if(bus_readOccur) begin
          mapping_claim_payload = targets_1_claim;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mapping_completion_valid = 1'b0;
    if(mapping_targetMapping_0_targetCompletion_valid) begin
      mapping_completion_valid = 1'b1;
    end
    if(mapping_targetMapping_1_targetCompletion_valid) begin
      mapping_completion_valid = 1'b1;
    end
  end

  always @(*) begin
    mapping_completion_payload = 5'bxxxxx;
    if(mapping_targetMapping_0_targetCompletion_valid) begin
      mapping_completion_payload = mapping_targetMapping_0_targetCompletion_payload;
    end
    if(mapping_targetMapping_1_targetCompletion_valid) begin
      mapping_completion_payload = mapping_targetMapping_1_targetCompletion_payload;
    end
  end

  always @(*) begin
    mapping_coherencyStall_willIncrement = 1'b0;
    if(when_PlicMapper_l122) begin
      mapping_coherencyStall_willIncrement = 1'b1;
    end
    if(when_AxiLite4SlaveFactory_l68) begin
      if(bus_writeJoinEvent_valid) begin
        mapping_coherencyStall_willIncrement = 1'b1;
      end
    end
    if(when_AxiLite4SlaveFactory_l86) begin
      if(bus_readDataStage_valid) begin
        mapping_coherencyStall_willIncrement = 1'b1;
      end
    end
  end

  assign mapping_coherencyStall_willClear = 1'b0;
  assign mapping_coherencyStall_willOverflowIfInc = (mapping_coherencyStall_value == 1'b1);
  assign mapping_coherencyStall_willOverflow = (mapping_coherencyStall_willOverflowIfInc && mapping_coherencyStall_willIncrement);
  always @(*) begin
    mapping_coherencyStall_valueNext = (mapping_coherencyStall_value + mapping_coherencyStall_willIncrement);
    if(mapping_coherencyStall_willClear) begin
      mapping_coherencyStall_valueNext = 1'b0;
    end
  end

  assign when_PlicMapper_l122 = (mapping_coherencyStall_value != 1'b0);
  assign targets_0_threshold = _zz_targets_0_threshold;
  always @(*) begin
    mapping_targetMapping_0_targetCompletion_valid = 1'b0;
    case(bus_writeAddressMasked)
      22'h200004 : begin
        if(bus_writeOccur) begin
          mapping_targetMapping_0_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign targets_0_ie_0 = _zz_targets_0_ie_0;
  assign targets_0_ie_1 = _zz_targets_0_ie_1;
  assign targets_0_ie_2 = _zz_targets_0_ie_2;
  assign targets_0_ie_3 = _zz_targets_0_ie_3;
  assign targets_0_ie_4 = _zz_targets_0_ie_4;
  assign targets_0_ie_5 = _zz_targets_0_ie_5;
  assign targets_0_ie_6 = _zz_targets_0_ie_6;
  assign targets_0_ie_7 = _zz_targets_0_ie_7;
  assign targets_0_ie_8 = _zz_targets_0_ie_8;
  assign targets_0_ie_9 = _zz_targets_0_ie_9;
  assign targets_0_ie_10 = _zz_targets_0_ie_10;
  assign targets_0_ie_11 = _zz_targets_0_ie_11;
  assign targets_0_ie_12 = _zz_targets_0_ie_12;
  assign targets_0_ie_13 = _zz_targets_0_ie_13;
  assign targets_0_ie_14 = _zz_targets_0_ie_14;
  assign targets_0_ie_15 = _zz_targets_0_ie_15;
  assign targets_0_ie_16 = _zz_targets_0_ie_16;
  assign targets_0_ie_17 = _zz_targets_0_ie_17;
  assign targets_0_ie_18 = _zz_targets_0_ie_18;
  assign targets_0_ie_19 = _zz_targets_0_ie_19;
  assign targets_0_ie_20 = _zz_targets_0_ie_20;
  assign targets_0_ie_21 = _zz_targets_0_ie_21;
  assign targets_0_ie_22 = _zz_targets_0_ie_22;
  assign targets_0_ie_23 = _zz_targets_0_ie_23;
  assign targets_0_ie_24 = _zz_targets_0_ie_24;
  assign targets_0_ie_25 = _zz_targets_0_ie_25;
  assign targets_0_ie_26 = _zz_targets_0_ie_26;
  assign targets_0_ie_27 = _zz_targets_0_ie_27;
  assign targets_0_ie_28 = _zz_targets_0_ie_28;
  assign targets_0_ie_29 = _zz_targets_0_ie_29;
  assign targets_0_ie_30 = _zz_targets_0_ie_30;
  assign targets_1_threshold = _zz_targets_1_threshold;
  always @(*) begin
    mapping_targetMapping_1_targetCompletion_valid = 1'b0;
    case(bus_writeAddressMasked)
      22'h201004 : begin
        if(bus_writeOccur) begin
          mapping_targetMapping_1_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign targets_1_ie_0 = _zz_targets_1_ie_0;
  assign targets_1_ie_1 = _zz_targets_1_ie_1;
  assign targets_1_ie_2 = _zz_targets_1_ie_2;
  assign targets_1_ie_3 = _zz_targets_1_ie_3;
  assign targets_1_ie_4 = _zz_targets_1_ie_4;
  assign targets_1_ie_5 = _zz_targets_1_ie_5;
  assign targets_1_ie_6 = _zz_targets_1_ie_6;
  assign targets_1_ie_7 = _zz_targets_1_ie_7;
  assign targets_1_ie_8 = _zz_targets_1_ie_8;
  assign targets_1_ie_9 = _zz_targets_1_ie_9;
  assign targets_1_ie_10 = _zz_targets_1_ie_10;
  assign targets_1_ie_11 = _zz_targets_1_ie_11;
  assign targets_1_ie_12 = _zz_targets_1_ie_12;
  assign targets_1_ie_13 = _zz_targets_1_ie_13;
  assign targets_1_ie_14 = _zz_targets_1_ie_14;
  assign targets_1_ie_15 = _zz_targets_1_ie_15;
  assign targets_1_ie_16 = _zz_targets_1_ie_16;
  assign targets_1_ie_17 = _zz_targets_1_ie_17;
  assign targets_1_ie_18 = _zz_targets_1_ie_18;
  assign targets_1_ie_19 = _zz_targets_1_ie_19;
  assign targets_1_ie_20 = _zz_targets_1_ie_20;
  assign targets_1_ie_21 = _zz_targets_1_ie_21;
  assign targets_1_ie_22 = _zz_targets_1_ie_22;
  assign targets_1_ie_23 = _zz_targets_1_ie_23;
  assign targets_1_ie_24 = _zz_targets_1_ie_24;
  assign targets_1_ie_25 = _zz_targets_1_ie_25;
  assign targets_1_ie_26 = _zz_targets_1_ie_26;
  assign targets_1_ie_27 = _zz_targets_1_ie_27;
  assign targets_1_ie_28 = _zz_targets_1_ie_28;
  assign targets_1_ie_29 = _zz_targets_1_ie_29;
  assign targets_1_ie_30 = _zz_targets_1_ie_30;
  assign mapping_targetMapping_0_targetCompletion_payload = io_bus_w_payload_data[4 : 0];
  assign mapping_targetMapping_1_targetCompletion_payload = io_bus_w_payload_data[4 : 0];
  assign when_AxiLite4SlaveFactory_l68 = 1'b1;
  assign when_AxiLite4SlaveFactory_l86 = 1'b1;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      gateways_0_ip <= 1'b0;
      gateways_0_waitCompletion <= 1'b0;
      gateways_1_ip <= 1'b0;
      gateways_1_waitCompletion <= 1'b0;
      gateways_2_ip <= 1'b0;
      gateways_2_waitCompletion <= 1'b0;
      gateways_3_ip <= 1'b0;
      gateways_3_waitCompletion <= 1'b0;
      gateways_4_ip <= 1'b0;
      gateways_4_waitCompletion <= 1'b0;
      gateways_5_ip <= 1'b0;
      gateways_5_waitCompletion <= 1'b0;
      gateways_6_ip <= 1'b0;
      gateways_6_waitCompletion <= 1'b0;
      gateways_7_ip <= 1'b0;
      gateways_7_waitCompletion <= 1'b0;
      gateways_8_ip <= 1'b0;
      gateways_8_waitCompletion <= 1'b0;
      gateways_9_ip <= 1'b0;
      gateways_9_waitCompletion <= 1'b0;
      gateways_10_ip <= 1'b0;
      gateways_10_waitCompletion <= 1'b0;
      gateways_11_ip <= 1'b0;
      gateways_11_waitCompletion <= 1'b0;
      gateways_12_ip <= 1'b0;
      gateways_12_waitCompletion <= 1'b0;
      gateways_13_ip <= 1'b0;
      gateways_13_waitCompletion <= 1'b0;
      gateways_14_ip <= 1'b0;
      gateways_14_waitCompletion <= 1'b0;
      gateways_15_ip <= 1'b0;
      gateways_15_waitCompletion <= 1'b0;
      gateways_16_ip <= 1'b0;
      gateways_16_waitCompletion <= 1'b0;
      gateways_17_ip <= 1'b0;
      gateways_17_waitCompletion <= 1'b0;
      gateways_18_ip <= 1'b0;
      gateways_18_waitCompletion <= 1'b0;
      gateways_19_ip <= 1'b0;
      gateways_19_waitCompletion <= 1'b0;
      gateways_20_ip <= 1'b0;
      gateways_20_waitCompletion <= 1'b0;
      gateways_21_ip <= 1'b0;
      gateways_21_waitCompletion <= 1'b0;
      gateways_22_ip <= 1'b0;
      gateways_22_waitCompletion <= 1'b0;
      gateways_23_ip <= 1'b0;
      gateways_23_waitCompletion <= 1'b0;
      gateways_24_ip <= 1'b0;
      gateways_24_waitCompletion <= 1'b0;
      gateways_25_ip <= 1'b0;
      gateways_25_waitCompletion <= 1'b0;
      gateways_26_ip <= 1'b0;
      gateways_26_waitCompletion <= 1'b0;
      gateways_27_ip <= 1'b0;
      gateways_27_waitCompletion <= 1'b0;
      gateways_28_ip <= 1'b0;
      gateways_28_waitCompletion <= 1'b0;
      gateways_29_ip <= 1'b0;
      gateways_29_waitCompletion <= 1'b0;
      gateways_30_ip <= 1'b0;
      gateways_30_waitCompletion <= 1'b0;
      _zz_io_bus_b_valid_1 <= 1'b0;
      io_bus_ar_rValid <= 1'b0;
      _zz_gateways_0_priority <= 2'b00;
      _zz_gateways_1_priority <= 2'b00;
      _zz_gateways_2_priority <= 2'b00;
      _zz_gateways_3_priority <= 2'b00;
      _zz_gateways_4_priority <= 2'b00;
      _zz_gateways_5_priority <= 2'b00;
      _zz_gateways_6_priority <= 2'b00;
      _zz_gateways_7_priority <= 2'b00;
      _zz_gateways_8_priority <= 2'b00;
      _zz_gateways_9_priority <= 2'b00;
      _zz_gateways_10_priority <= 2'b00;
      _zz_gateways_11_priority <= 2'b00;
      _zz_gateways_12_priority <= 2'b00;
      _zz_gateways_13_priority <= 2'b00;
      _zz_gateways_14_priority <= 2'b00;
      _zz_gateways_15_priority <= 2'b00;
      _zz_gateways_16_priority <= 2'b00;
      _zz_gateways_17_priority <= 2'b00;
      _zz_gateways_18_priority <= 2'b00;
      _zz_gateways_19_priority <= 2'b00;
      _zz_gateways_20_priority <= 2'b00;
      _zz_gateways_21_priority <= 2'b00;
      _zz_gateways_22_priority <= 2'b00;
      _zz_gateways_23_priority <= 2'b00;
      _zz_gateways_24_priority <= 2'b00;
      _zz_gateways_25_priority <= 2'b00;
      _zz_gateways_26_priority <= 2'b00;
      _zz_gateways_27_priority <= 2'b00;
      _zz_gateways_28_priority <= 2'b00;
      _zz_gateways_29_priority <= 2'b00;
      _zz_gateways_30_priority <= 2'b00;
      mapping_coherencyStall_value <= 1'b0;
      _zz_targets_0_threshold <= 2'b00;
      _zz_targets_0_ie_0 <= 1'b0;
      _zz_targets_0_ie_1 <= 1'b0;
      _zz_targets_0_ie_2 <= 1'b0;
      _zz_targets_0_ie_3 <= 1'b0;
      _zz_targets_0_ie_4 <= 1'b0;
      _zz_targets_0_ie_5 <= 1'b0;
      _zz_targets_0_ie_6 <= 1'b0;
      _zz_targets_0_ie_7 <= 1'b0;
      _zz_targets_0_ie_8 <= 1'b0;
      _zz_targets_0_ie_9 <= 1'b0;
      _zz_targets_0_ie_10 <= 1'b0;
      _zz_targets_0_ie_11 <= 1'b0;
      _zz_targets_0_ie_12 <= 1'b0;
      _zz_targets_0_ie_13 <= 1'b0;
      _zz_targets_0_ie_14 <= 1'b0;
      _zz_targets_0_ie_15 <= 1'b0;
      _zz_targets_0_ie_16 <= 1'b0;
      _zz_targets_0_ie_17 <= 1'b0;
      _zz_targets_0_ie_18 <= 1'b0;
      _zz_targets_0_ie_19 <= 1'b0;
      _zz_targets_0_ie_20 <= 1'b0;
      _zz_targets_0_ie_21 <= 1'b0;
      _zz_targets_0_ie_22 <= 1'b0;
      _zz_targets_0_ie_23 <= 1'b0;
      _zz_targets_0_ie_24 <= 1'b0;
      _zz_targets_0_ie_25 <= 1'b0;
      _zz_targets_0_ie_26 <= 1'b0;
      _zz_targets_0_ie_27 <= 1'b0;
      _zz_targets_0_ie_28 <= 1'b0;
      _zz_targets_0_ie_29 <= 1'b0;
      _zz_targets_0_ie_30 <= 1'b0;
      _zz_targets_1_threshold <= 2'b00;
      _zz_targets_1_ie_0 <= 1'b0;
      _zz_targets_1_ie_1 <= 1'b0;
      _zz_targets_1_ie_2 <= 1'b0;
      _zz_targets_1_ie_3 <= 1'b0;
      _zz_targets_1_ie_4 <= 1'b0;
      _zz_targets_1_ie_5 <= 1'b0;
      _zz_targets_1_ie_6 <= 1'b0;
      _zz_targets_1_ie_7 <= 1'b0;
      _zz_targets_1_ie_8 <= 1'b0;
      _zz_targets_1_ie_9 <= 1'b0;
      _zz_targets_1_ie_10 <= 1'b0;
      _zz_targets_1_ie_11 <= 1'b0;
      _zz_targets_1_ie_12 <= 1'b0;
      _zz_targets_1_ie_13 <= 1'b0;
      _zz_targets_1_ie_14 <= 1'b0;
      _zz_targets_1_ie_15 <= 1'b0;
      _zz_targets_1_ie_16 <= 1'b0;
      _zz_targets_1_ie_17 <= 1'b0;
      _zz_targets_1_ie_18 <= 1'b0;
      _zz_targets_1_ie_19 <= 1'b0;
      _zz_targets_1_ie_20 <= 1'b0;
      _zz_targets_1_ie_21 <= 1'b0;
      _zz_targets_1_ie_22 <= 1'b0;
      _zz_targets_1_ie_23 <= 1'b0;
      _zz_targets_1_ie_24 <= 1'b0;
      _zz_targets_1_ie_25 <= 1'b0;
      _zz_targets_1_ie_26 <= 1'b0;
      _zz_targets_1_ie_27 <= 1'b0;
      _zz_targets_1_ie_28 <= 1'b0;
      _zz_targets_1_ie_29 <= 1'b0;
      _zz_targets_1_ie_30 <= 1'b0;
    end else begin
      if(when_PlicGateway_l21) begin
        gateways_0_ip <= _zz_gateways_0_ip;
        gateways_0_waitCompletion <= _zz_gateways_0_ip;
      end
      if(when_PlicGateway_l21_1) begin
        gateways_1_ip <= _zz_gateways_1_ip;
        gateways_1_waitCompletion <= _zz_gateways_1_ip;
      end
      if(when_PlicGateway_l21_2) begin
        gateways_2_ip <= _zz_gateways_2_ip;
        gateways_2_waitCompletion <= _zz_gateways_2_ip;
      end
      if(when_PlicGateway_l21_3) begin
        gateways_3_ip <= _zz_gateways_3_ip;
        gateways_3_waitCompletion <= _zz_gateways_3_ip;
      end
      if(when_PlicGateway_l21_4) begin
        gateways_4_ip <= _zz_gateways_4_ip;
        gateways_4_waitCompletion <= _zz_gateways_4_ip;
      end
      if(when_PlicGateway_l21_5) begin
        gateways_5_ip <= _zz_gateways_5_ip;
        gateways_5_waitCompletion <= _zz_gateways_5_ip;
      end
      if(when_PlicGateway_l21_6) begin
        gateways_6_ip <= _zz_gateways_6_ip;
        gateways_6_waitCompletion <= _zz_gateways_6_ip;
      end
      if(when_PlicGateway_l21_7) begin
        gateways_7_ip <= _zz_gateways_7_ip;
        gateways_7_waitCompletion <= _zz_gateways_7_ip;
      end
      if(when_PlicGateway_l21_8) begin
        gateways_8_ip <= _zz_gateways_8_ip;
        gateways_8_waitCompletion <= _zz_gateways_8_ip;
      end
      if(when_PlicGateway_l21_9) begin
        gateways_9_ip <= _zz_gateways_9_ip;
        gateways_9_waitCompletion <= _zz_gateways_9_ip;
      end
      if(when_PlicGateway_l21_10) begin
        gateways_10_ip <= _zz_gateways_10_ip;
        gateways_10_waitCompletion <= _zz_gateways_10_ip;
      end
      if(when_PlicGateway_l21_11) begin
        gateways_11_ip <= _zz_gateways_11_ip;
        gateways_11_waitCompletion <= _zz_gateways_11_ip;
      end
      if(when_PlicGateway_l21_12) begin
        gateways_12_ip <= _zz_gateways_12_ip;
        gateways_12_waitCompletion <= _zz_gateways_12_ip;
      end
      if(when_PlicGateway_l21_13) begin
        gateways_13_ip <= _zz_gateways_13_ip;
        gateways_13_waitCompletion <= _zz_gateways_13_ip;
      end
      if(when_PlicGateway_l21_14) begin
        gateways_14_ip <= _zz_gateways_14_ip;
        gateways_14_waitCompletion <= _zz_gateways_14_ip;
      end
      if(when_PlicGateway_l21_15) begin
        gateways_15_ip <= _zz_gateways_15_ip;
        gateways_15_waitCompletion <= _zz_gateways_15_ip;
      end
      if(when_PlicGateway_l21_16) begin
        gateways_16_ip <= _zz_gateways_16_ip;
        gateways_16_waitCompletion <= _zz_gateways_16_ip;
      end
      if(when_PlicGateway_l21_17) begin
        gateways_17_ip <= _zz_gateways_17_ip;
        gateways_17_waitCompletion <= _zz_gateways_17_ip;
      end
      if(when_PlicGateway_l21_18) begin
        gateways_18_ip <= _zz_gateways_18_ip;
        gateways_18_waitCompletion <= _zz_gateways_18_ip;
      end
      if(when_PlicGateway_l21_19) begin
        gateways_19_ip <= _zz_gateways_19_ip;
        gateways_19_waitCompletion <= _zz_gateways_19_ip;
      end
      if(when_PlicGateway_l21_20) begin
        gateways_20_ip <= _zz_gateways_20_ip;
        gateways_20_waitCompletion <= _zz_gateways_20_ip;
      end
      if(when_PlicGateway_l21_21) begin
        gateways_21_ip <= _zz_gateways_21_ip;
        gateways_21_waitCompletion <= _zz_gateways_21_ip;
      end
      if(when_PlicGateway_l21_22) begin
        gateways_22_ip <= _zz_gateways_22_ip;
        gateways_22_waitCompletion <= _zz_gateways_22_ip;
      end
      if(when_PlicGateway_l21_23) begin
        gateways_23_ip <= _zz_gateways_23_ip;
        gateways_23_waitCompletion <= _zz_gateways_23_ip;
      end
      if(when_PlicGateway_l21_24) begin
        gateways_24_ip <= _zz_gateways_24_ip;
        gateways_24_waitCompletion <= _zz_gateways_24_ip;
      end
      if(when_PlicGateway_l21_25) begin
        gateways_25_ip <= _zz_gateways_25_ip;
        gateways_25_waitCompletion <= _zz_gateways_25_ip;
      end
      if(when_PlicGateway_l21_26) begin
        gateways_26_ip <= _zz_gateways_26_ip;
        gateways_26_waitCompletion <= _zz_gateways_26_ip;
      end
      if(when_PlicGateway_l21_27) begin
        gateways_27_ip <= _zz_gateways_27_ip;
        gateways_27_waitCompletion <= _zz_gateways_27_ip;
      end
      if(when_PlicGateway_l21_28) begin
        gateways_28_ip <= _zz_gateways_28_ip;
        gateways_28_waitCompletion <= _zz_gateways_28_ip;
      end
      if(when_PlicGateway_l21_29) begin
        gateways_29_ip <= _zz_gateways_29_ip;
        gateways_29_waitCompletion <= _zz_gateways_29_ip;
      end
      if(when_PlicGateway_l21_30) begin
        gateways_30_ip <= _zz_gateways_30_ip;
        gateways_30_waitCompletion <= _zz_gateways_30_ip;
      end
      if((bus_writeJoinEvent_translated_valid && _zz_bus_writeJoinEvent_translated_ready)) begin
        _zz_io_bus_b_valid_1 <= 1'b1;
      end
      if((_zz_io_bus_b_valid && io_bus_b_ready)) begin
        _zz_io_bus_b_valid_1 <= 1'b0;
      end
      if(io_bus_ar_valid) begin
        io_bus_ar_rValid <= 1'b1;
      end
      if(bus_readDataStage_fire) begin
        io_bus_ar_rValid <= 1'b0;
      end
      if(mapping_claim_valid) begin
        case(mapping_claim_payload)
          5'h01 : begin
            gateways_0_ip <= 1'b0;
          end
          5'h02 : begin
            gateways_1_ip <= 1'b0;
          end
          5'h03 : begin
            gateways_2_ip <= 1'b0;
          end
          5'h04 : begin
            gateways_3_ip <= 1'b0;
          end
          5'h05 : begin
            gateways_4_ip <= 1'b0;
          end
          5'h06 : begin
            gateways_5_ip <= 1'b0;
          end
          5'h07 : begin
            gateways_6_ip <= 1'b0;
          end
          5'h08 : begin
            gateways_7_ip <= 1'b0;
          end
          5'h09 : begin
            gateways_8_ip <= 1'b0;
          end
          5'h0a : begin
            gateways_9_ip <= 1'b0;
          end
          5'h0b : begin
            gateways_10_ip <= 1'b0;
          end
          5'h0c : begin
            gateways_11_ip <= 1'b0;
          end
          5'h0d : begin
            gateways_12_ip <= 1'b0;
          end
          5'h0e : begin
            gateways_13_ip <= 1'b0;
          end
          5'h0f : begin
            gateways_14_ip <= 1'b0;
          end
          5'h10 : begin
            gateways_15_ip <= 1'b0;
          end
          5'h11 : begin
            gateways_16_ip <= 1'b0;
          end
          5'h12 : begin
            gateways_17_ip <= 1'b0;
          end
          5'h13 : begin
            gateways_18_ip <= 1'b0;
          end
          5'h14 : begin
            gateways_19_ip <= 1'b0;
          end
          5'h15 : begin
            gateways_20_ip <= 1'b0;
          end
          5'h16 : begin
            gateways_21_ip <= 1'b0;
          end
          5'h17 : begin
            gateways_22_ip <= 1'b0;
          end
          5'h18 : begin
            gateways_23_ip <= 1'b0;
          end
          5'h19 : begin
            gateways_24_ip <= 1'b0;
          end
          5'h1a : begin
            gateways_25_ip <= 1'b0;
          end
          5'h1b : begin
            gateways_26_ip <= 1'b0;
          end
          5'h1c : begin
            gateways_27_ip <= 1'b0;
          end
          5'h1d : begin
            gateways_28_ip <= 1'b0;
          end
          5'h1e : begin
            gateways_29_ip <= 1'b0;
          end
          5'h1f : begin
            gateways_30_ip <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      if(mapping_completion_valid) begin
        case(mapping_completion_payload)
          5'h01 : begin
            gateways_0_waitCompletion <= 1'b0;
          end
          5'h02 : begin
            gateways_1_waitCompletion <= 1'b0;
          end
          5'h03 : begin
            gateways_2_waitCompletion <= 1'b0;
          end
          5'h04 : begin
            gateways_3_waitCompletion <= 1'b0;
          end
          5'h05 : begin
            gateways_4_waitCompletion <= 1'b0;
          end
          5'h06 : begin
            gateways_5_waitCompletion <= 1'b0;
          end
          5'h07 : begin
            gateways_6_waitCompletion <= 1'b0;
          end
          5'h08 : begin
            gateways_7_waitCompletion <= 1'b0;
          end
          5'h09 : begin
            gateways_8_waitCompletion <= 1'b0;
          end
          5'h0a : begin
            gateways_9_waitCompletion <= 1'b0;
          end
          5'h0b : begin
            gateways_10_waitCompletion <= 1'b0;
          end
          5'h0c : begin
            gateways_11_waitCompletion <= 1'b0;
          end
          5'h0d : begin
            gateways_12_waitCompletion <= 1'b0;
          end
          5'h0e : begin
            gateways_13_waitCompletion <= 1'b0;
          end
          5'h0f : begin
            gateways_14_waitCompletion <= 1'b0;
          end
          5'h10 : begin
            gateways_15_waitCompletion <= 1'b0;
          end
          5'h11 : begin
            gateways_16_waitCompletion <= 1'b0;
          end
          5'h12 : begin
            gateways_17_waitCompletion <= 1'b0;
          end
          5'h13 : begin
            gateways_18_waitCompletion <= 1'b0;
          end
          5'h14 : begin
            gateways_19_waitCompletion <= 1'b0;
          end
          5'h15 : begin
            gateways_20_waitCompletion <= 1'b0;
          end
          5'h16 : begin
            gateways_21_waitCompletion <= 1'b0;
          end
          5'h17 : begin
            gateways_22_waitCompletion <= 1'b0;
          end
          5'h18 : begin
            gateways_23_waitCompletion <= 1'b0;
          end
          5'h19 : begin
            gateways_24_waitCompletion <= 1'b0;
          end
          5'h1a : begin
            gateways_25_waitCompletion <= 1'b0;
          end
          5'h1b : begin
            gateways_26_waitCompletion <= 1'b0;
          end
          5'h1c : begin
            gateways_27_waitCompletion <= 1'b0;
          end
          5'h1d : begin
            gateways_28_waitCompletion <= 1'b0;
          end
          5'h1e : begin
            gateways_29_waitCompletion <= 1'b0;
          end
          5'h1f : begin
            gateways_30_waitCompletion <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      mapping_coherencyStall_value <= mapping_coherencyStall_valueNext;
      case(bus_writeAddressMasked)
        22'h000004 : begin
          if(bus_writeOccur) begin
            _zz_gateways_0_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000008 : begin
          if(bus_writeOccur) begin
            _zz_gateways_1_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h00000c : begin
          if(bus_writeOccur) begin
            _zz_gateways_2_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000010 : begin
          if(bus_writeOccur) begin
            _zz_gateways_3_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000014 : begin
          if(bus_writeOccur) begin
            _zz_gateways_4_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000018 : begin
          if(bus_writeOccur) begin
            _zz_gateways_5_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h00001c : begin
          if(bus_writeOccur) begin
            _zz_gateways_6_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000020 : begin
          if(bus_writeOccur) begin
            _zz_gateways_7_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000024 : begin
          if(bus_writeOccur) begin
            _zz_gateways_8_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000028 : begin
          if(bus_writeOccur) begin
            _zz_gateways_9_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h00002c : begin
          if(bus_writeOccur) begin
            _zz_gateways_10_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000030 : begin
          if(bus_writeOccur) begin
            _zz_gateways_11_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000034 : begin
          if(bus_writeOccur) begin
            _zz_gateways_12_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000038 : begin
          if(bus_writeOccur) begin
            _zz_gateways_13_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h00003c : begin
          if(bus_writeOccur) begin
            _zz_gateways_14_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000040 : begin
          if(bus_writeOccur) begin
            _zz_gateways_15_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000044 : begin
          if(bus_writeOccur) begin
            _zz_gateways_16_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000048 : begin
          if(bus_writeOccur) begin
            _zz_gateways_17_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h00004c : begin
          if(bus_writeOccur) begin
            _zz_gateways_18_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000050 : begin
          if(bus_writeOccur) begin
            _zz_gateways_19_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000054 : begin
          if(bus_writeOccur) begin
            _zz_gateways_20_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000058 : begin
          if(bus_writeOccur) begin
            _zz_gateways_21_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h00005c : begin
          if(bus_writeOccur) begin
            _zz_gateways_22_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000060 : begin
          if(bus_writeOccur) begin
            _zz_gateways_23_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000064 : begin
          if(bus_writeOccur) begin
            _zz_gateways_24_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000068 : begin
          if(bus_writeOccur) begin
            _zz_gateways_25_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h00006c : begin
          if(bus_writeOccur) begin
            _zz_gateways_26_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000070 : begin
          if(bus_writeOccur) begin
            _zz_gateways_27_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000074 : begin
          if(bus_writeOccur) begin
            _zz_gateways_28_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h000078 : begin
          if(bus_writeOccur) begin
            _zz_gateways_29_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h00007c : begin
          if(bus_writeOccur) begin
            _zz_gateways_30_priority <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h200000 : begin
          if(bus_writeOccur) begin
            _zz_targets_0_threshold <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h002000 : begin
          if(bus_writeOccur) begin
            _zz_targets_0_ie_0 <= io_bus_w_payload_data[1];
            _zz_targets_0_ie_1 <= io_bus_w_payload_data[2];
            _zz_targets_0_ie_2 <= io_bus_w_payload_data[3];
            _zz_targets_0_ie_3 <= io_bus_w_payload_data[4];
            _zz_targets_0_ie_4 <= io_bus_w_payload_data[5];
            _zz_targets_0_ie_5 <= io_bus_w_payload_data[6];
            _zz_targets_0_ie_6 <= io_bus_w_payload_data[7];
            _zz_targets_0_ie_7 <= io_bus_w_payload_data[8];
            _zz_targets_0_ie_8 <= io_bus_w_payload_data[9];
            _zz_targets_0_ie_9 <= io_bus_w_payload_data[10];
            _zz_targets_0_ie_10 <= io_bus_w_payload_data[11];
            _zz_targets_0_ie_11 <= io_bus_w_payload_data[12];
            _zz_targets_0_ie_12 <= io_bus_w_payload_data[13];
            _zz_targets_0_ie_13 <= io_bus_w_payload_data[14];
            _zz_targets_0_ie_14 <= io_bus_w_payload_data[15];
            _zz_targets_0_ie_15 <= io_bus_w_payload_data[16];
            _zz_targets_0_ie_16 <= io_bus_w_payload_data[17];
            _zz_targets_0_ie_17 <= io_bus_w_payload_data[18];
            _zz_targets_0_ie_18 <= io_bus_w_payload_data[19];
            _zz_targets_0_ie_19 <= io_bus_w_payload_data[20];
            _zz_targets_0_ie_20 <= io_bus_w_payload_data[21];
            _zz_targets_0_ie_21 <= io_bus_w_payload_data[22];
            _zz_targets_0_ie_22 <= io_bus_w_payload_data[23];
            _zz_targets_0_ie_23 <= io_bus_w_payload_data[24];
            _zz_targets_0_ie_24 <= io_bus_w_payload_data[25];
            _zz_targets_0_ie_25 <= io_bus_w_payload_data[26];
            _zz_targets_0_ie_26 <= io_bus_w_payload_data[27];
            _zz_targets_0_ie_27 <= io_bus_w_payload_data[28];
            _zz_targets_0_ie_28 <= io_bus_w_payload_data[29];
            _zz_targets_0_ie_29 <= io_bus_w_payload_data[30];
            _zz_targets_0_ie_30 <= io_bus_w_payload_data[31];
          end
        end
        22'h201000 : begin
          if(bus_writeOccur) begin
            _zz_targets_1_threshold <= io_bus_w_payload_data[1 : 0];
          end
        end
        22'h002080 : begin
          if(bus_writeOccur) begin
            _zz_targets_1_ie_0 <= io_bus_w_payload_data[1];
            _zz_targets_1_ie_1 <= io_bus_w_payload_data[2];
            _zz_targets_1_ie_2 <= io_bus_w_payload_data[3];
            _zz_targets_1_ie_3 <= io_bus_w_payload_data[4];
            _zz_targets_1_ie_4 <= io_bus_w_payload_data[5];
            _zz_targets_1_ie_5 <= io_bus_w_payload_data[6];
            _zz_targets_1_ie_6 <= io_bus_w_payload_data[7];
            _zz_targets_1_ie_7 <= io_bus_w_payload_data[8];
            _zz_targets_1_ie_8 <= io_bus_w_payload_data[9];
            _zz_targets_1_ie_9 <= io_bus_w_payload_data[10];
            _zz_targets_1_ie_10 <= io_bus_w_payload_data[11];
            _zz_targets_1_ie_11 <= io_bus_w_payload_data[12];
            _zz_targets_1_ie_12 <= io_bus_w_payload_data[13];
            _zz_targets_1_ie_13 <= io_bus_w_payload_data[14];
            _zz_targets_1_ie_14 <= io_bus_w_payload_data[15];
            _zz_targets_1_ie_15 <= io_bus_w_payload_data[16];
            _zz_targets_1_ie_16 <= io_bus_w_payload_data[17];
            _zz_targets_1_ie_17 <= io_bus_w_payload_data[18];
            _zz_targets_1_ie_18 <= io_bus_w_payload_data[19];
            _zz_targets_1_ie_19 <= io_bus_w_payload_data[20];
            _zz_targets_1_ie_20 <= io_bus_w_payload_data[21];
            _zz_targets_1_ie_21 <= io_bus_w_payload_data[22];
            _zz_targets_1_ie_22 <= io_bus_w_payload_data[23];
            _zz_targets_1_ie_23 <= io_bus_w_payload_data[24];
            _zz_targets_1_ie_24 <= io_bus_w_payload_data[25];
            _zz_targets_1_ie_25 <= io_bus_w_payload_data[26];
            _zz_targets_1_ie_26 <= io_bus_w_payload_data[27];
            _zz_targets_1_ie_27 <= io_bus_w_payload_data[28];
            _zz_targets_1_ie_28 <= io_bus_w_payload_data[29];
            _zz_targets_1_ie_29 <= io_bus_w_payload_data[30];
            _zz_targets_1_ie_30 <= io_bus_w_payload_data[31];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    targets_0_bestRequest_priority <= (_zz_targets_0_bestRequest_priority_6 ? _zz_targets_0_bestRequest_priority_4 : _zz_targets_0_bestRequest_priority_5);
    targets_0_bestRequest_id <= (_zz_targets_0_bestRequest_priority_6 ? (_zz_targets_0_bestRequest_id_80 ? (_zz_targets_0_bestRequest_id_72 ? (_zz_targets_0_bestRequest_id_48 ? _zz_targets_0_bestRequest_id_82 : _zz_targets_0_bestRequest_id_83) : (_zz_targets_0_bestRequest_id_51 ? _zz_targets_0_bestRequest_id_84 : _zz_targets_0_bestRequest_id_85)) : (_zz_targets_0_bestRequest_id_74 ? (_zz_targets_0_bestRequest_id_54 ? _zz_targets_0_bestRequest_id_86 : _zz_targets_0_bestRequest_id_87) : (_zz_targets_0_bestRequest_id_57 ? _zz_targets_0_bestRequest_id_88 : _zz_targets_0_bestRequest_id_89))) : (_zz_targets_0_bestRequest_id_81 ? (_zz_targets_0_bestRequest_id_76 ? (_zz_targets_0_bestRequest_id_60 ? _zz_targets_0_bestRequest_id_90 : _zz_targets_0_bestRequest_id_91) : (_zz_targets_0_bestRequest_id_63 ? _zz_targets_0_bestRequest_id_92 : _zz_targets_0_bestRequest_id_93)) : (_zz_targets_0_bestRequest_id_78 ? (_zz_targets_0_bestRequest_id_66 ? _zz_targets_0_bestRequest_id_94 : _zz_targets_0_bestRequest_id_95) : (_zz_targets_0_bestRequest_id_69 ? _zz_targets_0_bestRequest_id_96 : _zz_targets_0_bestRequest_id_97))));
    targets_0_bestRequest_valid <= (_zz_targets_0_bestRequest_priority_6 ? _zz_targets_0_bestRequest_valid : _zz_targets_0_bestRequest_valid_1);
    targets_1_bestRequest_priority <= (_zz_targets_1_bestRequest_priority_6 ? _zz_targets_1_bestRequest_priority_4 : _zz_targets_1_bestRequest_priority_5);
    targets_1_bestRequest_id <= (_zz_targets_1_bestRequest_priority_6 ? (_zz_targets_1_bestRequest_id_80 ? (_zz_targets_1_bestRequest_id_72 ? (_zz_targets_1_bestRequest_id_48 ? _zz_targets_1_bestRequest_id_82 : _zz_targets_1_bestRequest_id_83) : (_zz_targets_1_bestRequest_id_51 ? _zz_targets_1_bestRequest_id_84 : _zz_targets_1_bestRequest_id_85)) : (_zz_targets_1_bestRequest_id_74 ? (_zz_targets_1_bestRequest_id_54 ? _zz_targets_1_bestRequest_id_86 : _zz_targets_1_bestRequest_id_87) : (_zz_targets_1_bestRequest_id_57 ? _zz_targets_1_bestRequest_id_88 : _zz_targets_1_bestRequest_id_89))) : (_zz_targets_1_bestRequest_id_81 ? (_zz_targets_1_bestRequest_id_76 ? (_zz_targets_1_bestRequest_id_60 ? _zz_targets_1_bestRequest_id_90 : _zz_targets_1_bestRequest_id_91) : (_zz_targets_1_bestRequest_id_63 ? _zz_targets_1_bestRequest_id_92 : _zz_targets_1_bestRequest_id_93)) : (_zz_targets_1_bestRequest_id_78 ? (_zz_targets_1_bestRequest_id_66 ? _zz_targets_1_bestRequest_id_94 : _zz_targets_1_bestRequest_id_95) : (_zz_targets_1_bestRequest_id_69 ? _zz_targets_1_bestRequest_id_96 : _zz_targets_1_bestRequest_id_97))));
    targets_1_bestRequest_valid <= (_zz_targets_1_bestRequest_priority_6 ? _zz_targets_1_bestRequest_valid : _zz_targets_1_bestRequest_valid_1);
    if(_zz_bus_writeJoinEvent_translated_ready_1) begin
      _zz_io_bus_b_payload_resp <= bus_writeJoinEvent_translated_payload_resp;
    end
    if(io_bus_ar_ready) begin
      io_bus_ar_rData_addr <= io_bus_ar_payload_addr;
      io_bus_ar_rData_prot <= io_bus_ar_payload_prot;
    end
  end


endmodule

module AxiLite4Clint (
  input  wire          io_bus_aw_valid,
  output wire          io_bus_aw_ready,
  input  wire [15:0]   io_bus_aw_payload_addr,
  input  wire [2:0]    io_bus_aw_payload_prot,
  input  wire          io_bus_w_valid,
  output wire          io_bus_w_ready,
  input  wire [31:0]   io_bus_w_payload_data,
  input  wire [3:0]    io_bus_w_payload_strb,
  output wire          io_bus_b_valid,
  input  wire          io_bus_b_ready,
  output wire [1:0]    io_bus_b_payload_resp,
  input  wire          io_bus_ar_valid,
  output wire          io_bus_ar_ready,
  input  wire [15:0]   io_bus_ar_payload_addr,
  input  wire [2:0]    io_bus_ar_payload_prot,
  output wire          io_bus_r_valid,
  input  wire          io_bus_r_ready,
  output wire [31:0]   io_bus_r_payload_data,
  output wire [1:0]    io_bus_r_payload_resp,
  output wire [0:0]    io_timerInterrupt,
  output wire [0:0]    io_softwareInterrupt,
  output wire [63:0]   io_time,
  input  wire          clk,
  input  wire          reset
);

  wire                factory_readErrorFlag;
  wire                factory_writeErrorFlag;
  wire                factory_readHaltRequest;
  wire                factory_writeHaltRequest;
  wire                factory_writeJoinEvent_valid;
  wire                factory_writeJoinEvent_ready;
  wire                factory_writeOccur;
  reg        [1:0]    factory_writeRsp_resp;
  wire                factory_writeJoinEvent_translated_valid;
  wire                factory_writeJoinEvent_translated_ready;
  wire       [1:0]    factory_writeJoinEvent_translated_payload_resp;
  wire                _zz_factory_writeJoinEvent_translated_ready;
  wire                _zz_factory_writeJoinEvent_translated_ready_1;
  wire                _zz_io_bus_b_valid;
  reg                 _zz_io_bus_b_valid_1;
  reg        [1:0]    _zz_io_bus_b_payload_resp;
  wire                factory_readDataStage_valid;
  wire                factory_readDataStage_ready;
  wire       [15:0]   factory_readDataStage_payload_addr;
  wire       [2:0]    factory_readDataStage_payload_prot;
  reg                 io_bus_ar_rValid;
  wire                factory_readDataStage_fire;
  reg        [15:0]   io_bus_ar_rData_addr;
  reg        [2:0]    io_bus_ar_rData_prot;
  reg        [31:0]   factory_readRsp_data;
  reg        [1:0]    factory_readRsp_resp;
  wire                _zz_io_bus_r_valid;
  wire       [15:0]   factory_readAddressMasked;
  wire       [15:0]   factory_writeAddressMasked;
  wire                factory_readOccur;
  wire                logic_stop;
  reg        [63:0]   logic_time;
  wire                when_Clint_l39;
  reg        [63:0]   logic_harts_0_cmp;
  reg                 logic_harts_0_timerInterrupt;
  reg                 logic_harts_0_softwareInterrupt;
  wire       [63:0]   _zz_factory_readRsp_data;
  wire                when_AxiLite4SlaveFactory_l68;
  wire                when_AxiLite4SlaveFactory_l68_1;
  wire                when_AxiLite4SlaveFactory_l86;
  wire                when_AxiLite4SlaveFactory_l86_1;

  assign factory_readErrorFlag = 1'b0;
  assign factory_writeErrorFlag = 1'b0;
  assign factory_readHaltRequest = 1'b0;
  assign factory_writeHaltRequest = 1'b0;
  assign factory_writeOccur = (factory_writeJoinEvent_valid && factory_writeJoinEvent_ready);
  assign factory_writeJoinEvent_valid = (io_bus_aw_valid && io_bus_w_valid);
  assign io_bus_aw_ready = factory_writeOccur;
  assign io_bus_w_ready = factory_writeOccur;
  assign factory_writeJoinEvent_translated_valid = factory_writeJoinEvent_valid;
  assign factory_writeJoinEvent_ready = factory_writeJoinEvent_translated_ready;
  assign factory_writeJoinEvent_translated_payload_resp = factory_writeRsp_resp;
  assign _zz_factory_writeJoinEvent_translated_ready = (! factory_writeHaltRequest);
  assign factory_writeJoinEvent_translated_ready = (_zz_factory_writeJoinEvent_translated_ready_1 && _zz_factory_writeJoinEvent_translated_ready);
  assign _zz_factory_writeJoinEvent_translated_ready_1 = (! _zz_io_bus_b_valid_1);
  assign _zz_io_bus_b_valid = _zz_io_bus_b_valid_1;
  assign io_bus_b_valid = _zz_io_bus_b_valid;
  assign io_bus_b_payload_resp = _zz_io_bus_b_payload_resp;
  assign factory_readDataStage_fire = (factory_readDataStage_valid && factory_readDataStage_ready);
  assign io_bus_ar_ready = (! io_bus_ar_rValid);
  assign factory_readDataStage_valid = io_bus_ar_rValid;
  assign factory_readDataStage_payload_addr = io_bus_ar_rData_addr;
  assign factory_readDataStage_payload_prot = io_bus_ar_rData_prot;
  assign _zz_io_bus_r_valid = (! factory_readHaltRequest);
  assign factory_readDataStage_ready = (io_bus_r_ready && _zz_io_bus_r_valid);
  assign io_bus_r_valid = (factory_readDataStage_valid && _zz_io_bus_r_valid);
  assign io_bus_r_payload_data = factory_readRsp_data;
  assign io_bus_r_payload_resp = factory_readRsp_resp;
  always @(*) begin
    if(factory_writeErrorFlag) begin
      factory_writeRsp_resp = 2'b10;
    end else begin
      factory_writeRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    if(factory_readErrorFlag) begin
      factory_readRsp_resp = 2'b10;
    end else begin
      factory_readRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    factory_readRsp_data = 32'h00000000;
    case(factory_readAddressMasked)
      16'h0000 : begin
        factory_readRsp_data[0 : 0] = logic_harts_0_softwareInterrupt;
      end
      default : begin
      end
    endcase
    if(when_AxiLite4SlaveFactory_l86) begin
      factory_readRsp_data[31 : 0] = _zz_factory_readRsp_data[31 : 0];
    end
    if(when_AxiLite4SlaveFactory_l86_1) begin
      factory_readRsp_data[31 : 0] = _zz_factory_readRsp_data[63 : 32];
    end
  end

  assign factory_readAddressMasked = (factory_readDataStage_payload_addr & (~ 16'h0003));
  assign factory_writeAddressMasked = (io_bus_aw_payload_addr & (~ 16'h0003));
  assign factory_readOccur = (io_bus_r_valid && io_bus_r_ready);
  assign logic_stop = 1'b0;
  assign when_Clint_l39 = (! logic_stop);
  assign _zz_factory_readRsp_data = logic_time;
  assign io_timerInterrupt[0] = logic_harts_0_timerInterrupt;
  assign io_softwareInterrupt[0] = logic_harts_0_softwareInterrupt;
  assign io_time = logic_time;
  assign when_AxiLite4SlaveFactory_l68 = ((factory_writeAddressMasked & (~ 16'h0003)) == 16'h4000);
  assign when_AxiLite4SlaveFactory_l68_1 = ((factory_writeAddressMasked & (~ 16'h0003)) == 16'h4004);
  assign when_AxiLite4SlaveFactory_l86 = ((factory_readAddressMasked & (~ 16'h0003)) == 16'hbff8);
  assign when_AxiLite4SlaveFactory_l86_1 = ((factory_readAddressMasked & (~ 16'h0003)) == 16'hbffc);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _zz_io_bus_b_valid_1 <= 1'b0;
      io_bus_ar_rValid <= 1'b0;
      logic_time <= 64'h0000000000000000;
      logic_harts_0_softwareInterrupt <= 1'b0;
    end else begin
      if((factory_writeJoinEvent_translated_valid && _zz_factory_writeJoinEvent_translated_ready)) begin
        _zz_io_bus_b_valid_1 <= 1'b1;
      end
      if((_zz_io_bus_b_valid && io_bus_b_ready)) begin
        _zz_io_bus_b_valid_1 <= 1'b0;
      end
      if(io_bus_ar_valid) begin
        io_bus_ar_rValid <= 1'b1;
      end
      if(factory_readDataStage_fire) begin
        io_bus_ar_rValid <= 1'b0;
      end
      if(when_Clint_l39) begin
        logic_time <= (logic_time + 64'h0000000000000001);
      end
      case(factory_writeAddressMasked)
        16'h0000 : begin
          if(factory_writeOccur) begin
            logic_harts_0_softwareInterrupt <= io_bus_w_payload_data[0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if(_zz_factory_writeJoinEvent_translated_ready_1) begin
      _zz_io_bus_b_payload_resp <= factory_writeJoinEvent_translated_payload_resp;
    end
    if(io_bus_ar_ready) begin
      io_bus_ar_rData_addr <= io_bus_ar_payload_addr;
      io_bus_ar_rData_prot <= io_bus_ar_payload_prot;
    end
    logic_harts_0_timerInterrupt <= (logic_harts_0_cmp <= logic_time);
    if(when_AxiLite4SlaveFactory_l68) begin
      if(factory_writeOccur) begin
        logic_harts_0_cmp[31 : 0] <= io_bus_w_payload_data[31 : 0];
      end
    end
    if(when_AxiLite4SlaveFactory_l68_1) begin
      if(factory_writeOccur) begin
        logic_harts_0_cmp[63 : 32] <= io_bus_w_payload_data[31 : 0];
      end
    end
  end


endmodule

module StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [3:0]    io_push_payload_robId,
  input  wire [0:0]    io_push_payload_mask,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [3:0]    io_pop_payload_robId,
  output wire [0:0]    io_pop_payload_mask,
  input  wire          io_flush,
  output wire [4:0]    io_occupancy,
  output wire [4:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire       [4:0]    logic_ram_spinal_port1;
  wire       [4:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [4:0]    logic_ptr_push;
  reg        [4:0]    logic_ptr_pop;
  wire       [4:0]    logic_ptr_occupancy;
  wire       [4:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1243;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [3:0]    logic_push_onRam_write_payload_address;
  wire       [3:0]    logic_push_onRam_write_payload_data_robId;
  wire       [0:0]    logic_push_onRam_write_payload_data_mask;
  wire                logic_pop_addressGen_valid;
  wire                logic_pop_addressGen_ready;
  wire       [3:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire       [3:0]    logic_pop_async_readed_robId;
  wire       [0:0]    logic_pop_async_readed_mask;
  wire       [4:0]    _zz_logic_pop_async_readed_robId;
  wire                logic_pop_addressGen_translated_valid;
  wire                logic_pop_addressGen_translated_ready;
  wire       [3:0]    logic_pop_addressGen_translated_payload_robId;
  wire       [0:0]    logic_pop_addressGen_translated_payload_mask;
  (* ram_style = "distributed" *) reg [4:0] logic_ram [0:15];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_mask,logic_push_onRam_write_payload_data_robId};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  assign logic_ram_spinal_port1 = logic_ram[logic_pop_addressGen_payload];
  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1243 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 5'h10) == 5'h00);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[3:0];
  assign logic_push_onRam_write_payload_data_robId = io_push_payload_robId;
  assign logic_push_onRam_write_payload_data_mask = io_push_payload_mask;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[3:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  assign _zz_logic_pop_async_readed_robId = logic_ram_spinal_port1;
  assign logic_pop_async_readed_robId = _zz_logic_pop_async_readed_robId[3 : 0];
  assign logic_pop_async_readed_mask = _zz_logic_pop_async_readed_robId[4 : 4];
  assign logic_pop_addressGen_translated_valid = logic_pop_addressGen_valid;
  assign logic_pop_addressGen_ready = logic_pop_addressGen_translated_ready;
  assign logic_pop_addressGen_translated_payload_robId = logic_pop_async_readed_robId;
  assign logic_pop_addressGen_translated_payload_mask = logic_pop_async_readed_mask;
  assign io_pop_valid = logic_pop_addressGen_translated_valid;
  assign logic_pop_addressGen_translated_ready = io_pop_ready;
  assign io_pop_payload_robId = logic_pop_addressGen_translated_payload_robId;
  assign io_pop_payload_mask = logic_pop_addressGen_translated_payload_mask;
  assign logic_ptr_popOnIo = logic_ptr_pop;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (5'h10 - logic_ptr_occupancy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_ptr_push <= 5'h00;
      logic_ptr_pop <= 5'h00;
      logic_ptr_wentUp <= 1'b0;
    end else begin
      if(when_Stream_l1243) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 5'h01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 5'h01);
      end
      if(io_flush) begin
        logic_ptr_push <= 5'h00;
        logic_ptr_pop <= 5'h00;
      end
    end
  end


endmodule
